VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Proc
  CLASS BLOCK ;
  FOREIGN Proc ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.750 596.000 10.030 600.000 ;
    END
  END clk
  PIN dmemreq_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END dmemreq_addr[0]
  PIN dmemreq_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END dmemreq_addr[10]
  PIN dmemreq_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END dmemreq_addr[11]
  PIN dmemreq_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END dmemreq_addr[12]
  PIN dmemreq_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END dmemreq_addr[13]
  PIN dmemreq_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END dmemreq_addr[14]
  PIN dmemreq_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END dmemreq_addr[15]
  PIN dmemreq_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END dmemreq_addr[16]
  PIN dmemreq_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END dmemreq_addr[17]
  PIN dmemreq_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END dmemreq_addr[18]
  PIN dmemreq_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END dmemreq_addr[19]
  PIN dmemreq_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END dmemreq_addr[1]
  PIN dmemreq_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END dmemreq_addr[20]
  PIN dmemreq_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END dmemreq_addr[21]
  PIN dmemreq_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END dmemreq_addr[22]
  PIN dmemreq_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END dmemreq_addr[23]
  PIN dmemreq_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END dmemreq_addr[24]
  PIN dmemreq_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END dmemreq_addr[25]
  PIN dmemreq_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END dmemreq_addr[26]
  PIN dmemreq_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END dmemreq_addr[27]
  PIN dmemreq_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END dmemreq_addr[28]
  PIN dmemreq_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END dmemreq_addr[29]
  PIN dmemreq_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END dmemreq_addr[2]
  PIN dmemreq_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END dmemreq_addr[30]
  PIN dmemreq_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END dmemreq_addr[31]
  PIN dmemreq_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END dmemreq_addr[3]
  PIN dmemreq_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END dmemreq_addr[4]
  PIN dmemreq_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END dmemreq_addr[5]
  PIN dmemreq_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END dmemreq_addr[6]
  PIN dmemreq_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END dmemreq_addr[7]
  PIN dmemreq_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END dmemreq_addr[8]
  PIN dmemreq_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END dmemreq_addr[9]
  PIN dmemreq_type
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END dmemreq_type
  PIN dmemreq_val
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END dmemreq_val
  PIN dmemreq_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END dmemreq_wdata[0]
  PIN dmemreq_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END dmemreq_wdata[10]
  PIN dmemreq_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END dmemreq_wdata[11]
  PIN dmemreq_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END dmemreq_wdata[12]
  PIN dmemreq_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END dmemreq_wdata[13]
  PIN dmemreq_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END dmemreq_wdata[14]
  PIN dmemreq_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END dmemreq_wdata[15]
  PIN dmemreq_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END dmemreq_wdata[16]
  PIN dmemreq_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END dmemreq_wdata[17]
  PIN dmemreq_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END dmemreq_wdata[18]
  PIN dmemreq_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END dmemreq_wdata[19]
  PIN dmemreq_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END dmemreq_wdata[1]
  PIN dmemreq_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END dmemreq_wdata[20]
  PIN dmemreq_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END dmemreq_wdata[21]
  PIN dmemreq_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END dmemreq_wdata[22]
  PIN dmemreq_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END dmemreq_wdata[23]
  PIN dmemreq_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END dmemreq_wdata[24]
  PIN dmemreq_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END dmemreq_wdata[25]
  PIN dmemreq_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END dmemreq_wdata[26]
  PIN dmemreq_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END dmemreq_wdata[27]
  PIN dmemreq_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END dmemreq_wdata[28]
  PIN dmemreq_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END dmemreq_wdata[29]
  PIN dmemreq_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END dmemreq_wdata[2]
  PIN dmemreq_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END dmemreq_wdata[30]
  PIN dmemreq_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END dmemreq_wdata[31]
  PIN dmemreq_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END dmemreq_wdata[3]
  PIN dmemreq_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END dmemreq_wdata[4]
  PIN dmemreq_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END dmemreq_wdata[5]
  PIN dmemreq_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END dmemreq_wdata[6]
  PIN dmemreq_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END dmemreq_wdata[7]
  PIN dmemreq_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END dmemreq_wdata[8]
  PIN dmemreq_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END dmemreq_wdata[9]
  PIN dmemresp_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END dmemresp_rdata[0]
  PIN dmemresp_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END dmemresp_rdata[10]
  PIN dmemresp_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END dmemresp_rdata[11]
  PIN dmemresp_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END dmemresp_rdata[12]
  PIN dmemresp_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END dmemresp_rdata[13]
  PIN dmemresp_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END dmemresp_rdata[14]
  PIN dmemresp_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END dmemresp_rdata[15]
  PIN dmemresp_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END dmemresp_rdata[16]
  PIN dmemresp_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END dmemresp_rdata[17]
  PIN dmemresp_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END dmemresp_rdata[18]
  PIN dmemresp_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END dmemresp_rdata[19]
  PIN dmemresp_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END dmemresp_rdata[1]
  PIN dmemresp_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END dmemresp_rdata[20]
  PIN dmemresp_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END dmemresp_rdata[21]
  PIN dmemresp_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END dmemresp_rdata[22]
  PIN dmemresp_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END dmemresp_rdata[23]
  PIN dmemresp_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END dmemresp_rdata[24]
  PIN dmemresp_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END dmemresp_rdata[25]
  PIN dmemresp_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END dmemresp_rdata[26]
  PIN dmemresp_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END dmemresp_rdata[27]
  PIN dmemresp_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END dmemresp_rdata[28]
  PIN dmemresp_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END dmemresp_rdata[29]
  PIN dmemresp_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END dmemresp_rdata[2]
  PIN dmemresp_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END dmemresp_rdata[30]
  PIN dmemresp_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END dmemresp_rdata[31]
  PIN dmemresp_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END dmemresp_rdata[3]
  PIN dmemresp_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END dmemresp_rdata[4]
  PIN dmemresp_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END dmemresp_rdata[5]
  PIN dmemresp_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END dmemresp_rdata[6]
  PIN dmemresp_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END dmemresp_rdata[7]
  PIN dmemresp_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END dmemresp_rdata[8]
  PIN dmemresp_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END dmemresp_rdata[9]
  PIN imemreq_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END imemreq_addr[0]
  PIN imemreq_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END imemreq_addr[10]
  PIN imemreq_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END imemreq_addr[11]
  PIN imemreq_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END imemreq_addr[12]
  PIN imemreq_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END imemreq_addr[13]
  PIN imemreq_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END imemreq_addr[14]
  PIN imemreq_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END imemreq_addr[15]
  PIN imemreq_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END imemreq_addr[16]
  PIN imemreq_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END imemreq_addr[17]
  PIN imemreq_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END imemreq_addr[18]
  PIN imemreq_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END imemreq_addr[19]
  PIN imemreq_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END imemreq_addr[1]
  PIN imemreq_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END imemreq_addr[20]
  PIN imemreq_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END imemreq_addr[21]
  PIN imemreq_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END imemreq_addr[22]
  PIN imemreq_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END imemreq_addr[23]
  PIN imemreq_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END imemreq_addr[24]
  PIN imemreq_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END imemreq_addr[25]
  PIN imemreq_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END imemreq_addr[26]
  PIN imemreq_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END imemreq_addr[27]
  PIN imemreq_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END imemreq_addr[28]
  PIN imemreq_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END imemreq_addr[29]
  PIN imemreq_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END imemreq_addr[2]
  PIN imemreq_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END imemreq_addr[30]
  PIN imemreq_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END imemreq_addr[31]
  PIN imemreq_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END imemreq_addr[3]
  PIN imemreq_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END imemreq_addr[4]
  PIN imemreq_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END imemreq_addr[5]
  PIN imemreq_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END imemreq_addr[6]
  PIN imemreq_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END imemreq_addr[7]
  PIN imemreq_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END imemreq_addr[8]
  PIN imemreq_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END imemreq_addr[9]
  PIN imemreq_val
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END imemreq_val
  PIN imemresp_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END imemresp_data[0]
  PIN imemresp_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END imemresp_data[10]
  PIN imemresp_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END imemresp_data[11]
  PIN imemresp_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END imemresp_data[12]
  PIN imemresp_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END imemresp_data[13]
  PIN imemresp_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END imemresp_data[14]
  PIN imemresp_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END imemresp_data[15]
  PIN imemresp_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END imemresp_data[16]
  PIN imemresp_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END imemresp_data[17]
  PIN imemresp_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END imemresp_data[18]
  PIN imemresp_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END imemresp_data[19]
  PIN imemresp_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END imemresp_data[1]
  PIN imemresp_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END imemresp_data[20]
  PIN imemresp_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END imemresp_data[21]
  PIN imemresp_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END imemresp_data[22]
  PIN imemresp_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END imemresp_data[23]
  PIN imemresp_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END imemresp_data[24]
  PIN imemresp_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END imemresp_data[25]
  PIN imemresp_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END imemresp_data[26]
  PIN imemresp_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END imemresp_data[27]
  PIN imemresp_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END imemresp_data[28]
  PIN imemresp_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END imemresp_data[29]
  PIN imemresp_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END imemresp_data[2]
  PIN imemresp_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END imemresp_data[30]
  PIN imemresp_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END imemresp_data[31]
  PIN imemresp_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END imemresp_data[3]
  PIN imemresp_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END imemresp_data[4]
  PIN imemresp_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END imemresp_data[5]
  PIN imemresp_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END imemresp_data[6]
  PIN imemresp_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END imemresp_data[7]
  PIN imemresp_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END imemresp_data[8]
  PIN imemresp_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END imemresp_data[9]
  PIN in0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 21.710 596.000 21.990 600.000 ;
    END
  END in0[0]
  PIN in0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 596.000 81.790 600.000 ;
    END
  END in0[10]
  PIN in0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.490 596.000 87.770 600.000 ;
    END
  END in0[11]
  PIN in0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 596.000 93.750 600.000 ;
    END
  END in0[12]
  PIN in0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 596.000 99.730 600.000 ;
    END
  END in0[13]
  PIN in0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 105.430 596.000 105.710 600.000 ;
    END
  END in0[14]
  PIN in0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 596.000 111.690 600.000 ;
    END
  END in0[15]
  PIN in0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 117.390 596.000 117.670 600.000 ;
    END
  END in0[16]
  PIN in0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 123.370 596.000 123.650 600.000 ;
    END
  END in0[17]
  PIN in0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 129.350 596.000 129.630 600.000 ;
    END
  END in0[18]
  PIN in0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 596.000 135.610 600.000 ;
    END
  END in0[19]
  PIN in0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.690 596.000 27.970 600.000 ;
    END
  END in0[1]
  PIN in0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 141.310 596.000 141.590 600.000 ;
    END
  END in0[20]
  PIN in0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 147.290 596.000 147.570 600.000 ;
    END
  END in0[21]
  PIN in0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 596.000 153.550 600.000 ;
    END
  END in0[22]
  PIN in0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 596.000 159.530 600.000 ;
    END
  END in0[23]
  PIN in0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.230 596.000 165.510 600.000 ;
    END
  END in0[24]
  PIN in0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 171.210 596.000 171.490 600.000 ;
    END
  END in0[25]
  PIN in0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 596.000 177.470 600.000 ;
    END
  END in0[26]
  PIN in0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.170 596.000 183.450 600.000 ;
    END
  END in0[27]
  PIN in0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 189.150 596.000 189.430 600.000 ;
    END
  END in0[28]
  PIN in0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 596.000 195.410 600.000 ;
    END
  END in0[29]
  PIN in0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 596.000 33.950 600.000 ;
    END
  END in0[2]
  PIN in0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 201.110 596.000 201.390 600.000 ;
    END
  END in0[30]
  PIN in0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 207.090 596.000 207.370 600.000 ;
    END
  END in0[31]
  PIN in0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 596.000 39.930 600.000 ;
    END
  END in0[3]
  PIN in0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.630 596.000 45.910 600.000 ;
    END
  END in0[4]
  PIN in0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 596.000 51.890 600.000 ;
    END
  END in0[5]
  PIN in0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 57.590 596.000 57.870 600.000 ;
    END
  END in0[6]
  PIN in0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.570 596.000 63.850 600.000 ;
    END
  END in0[7]
  PIN in0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 69.550 596.000 69.830 600.000 ;
    END
  END in0[8]
  PIN in0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.530 596.000 75.810 600.000 ;
    END
  END in0[9]
  PIN in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 213.070 596.000 213.350 600.000 ;
    END
  END in1[0]
  PIN in1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 272.870 596.000 273.150 600.000 ;
    END
  END in1[10]
  PIN in1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 278.850 596.000 279.130 600.000 ;
    END
  END in1[11]
  PIN in1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 284.830 596.000 285.110 600.000 ;
    END
  END in1[12]
  PIN in1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 290.810 596.000 291.090 600.000 ;
    END
  END in1[13]
  PIN in1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 296.790 596.000 297.070 600.000 ;
    END
  END in1[14]
  PIN in1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 596.000 303.050 600.000 ;
    END
  END in1[15]
  PIN in1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 308.750 596.000 309.030 600.000 ;
    END
  END in1[16]
  PIN in1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 314.730 596.000 315.010 600.000 ;
    END
  END in1[17]
  PIN in1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 320.710 596.000 320.990 600.000 ;
    END
  END in1[18]
  PIN in1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 326.690 596.000 326.970 600.000 ;
    END
  END in1[19]
  PIN in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 596.000 219.330 600.000 ;
    END
  END in1[1]
  PIN in1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 332.670 596.000 332.950 600.000 ;
    END
  END in1[20]
  PIN in1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 338.650 596.000 338.930 600.000 ;
    END
  END in1[21]
  PIN in1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 344.630 596.000 344.910 600.000 ;
    END
  END in1[22]
  PIN in1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 350.610 596.000 350.890 600.000 ;
    END
  END in1[23]
  PIN in1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 356.590 596.000 356.870 600.000 ;
    END
  END in1[24]
  PIN in1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 362.570 596.000 362.850 600.000 ;
    END
  END in1[25]
  PIN in1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 368.550 596.000 368.830 600.000 ;
    END
  END in1[26]
  PIN in1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 374.530 596.000 374.810 600.000 ;
    END
  END in1[27]
  PIN in1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 380.510 596.000 380.790 600.000 ;
    END
  END in1[28]
  PIN in1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 596.000 386.770 600.000 ;
    END
  END in1[29]
  PIN in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.030 596.000 225.310 600.000 ;
    END
  END in1[2]
  PIN in1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 392.470 596.000 392.750 600.000 ;
    END
  END in1[30]
  PIN in1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 398.450 596.000 398.730 600.000 ;
    END
  END in1[31]
  PIN in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 231.010 596.000 231.290 600.000 ;
    END
  END in1[3]
  PIN in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 236.990 596.000 237.270 600.000 ;
    END
  END in1[4]
  PIN in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 242.970 596.000 243.250 600.000 ;
    END
  END in1[5]
  PIN in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.950 596.000 249.230 600.000 ;
    END
  END in1[6]
  PIN in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 254.930 596.000 255.210 600.000 ;
    END
  END in1[7]
  PIN in1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 260.910 596.000 261.190 600.000 ;
    END
  END in1[8]
  PIN in1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 266.890 596.000 267.170 600.000 ;
    END
  END in1[9]
  PIN in2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 404.430 596.000 404.710 600.000 ;
    END
  END in2[0]
  PIN in2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 464.230 596.000 464.510 600.000 ;
    END
  END in2[10]
  PIN in2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 596.000 470.490 600.000 ;
    END
  END in2[11]
  PIN in2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 476.190 596.000 476.470 600.000 ;
    END
  END in2[12]
  PIN in2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 596.000 482.450 600.000 ;
    END
  END in2[13]
  PIN in2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 488.150 596.000 488.430 600.000 ;
    END
  END in2[14]
  PIN in2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 596.000 494.410 600.000 ;
    END
  END in2[15]
  PIN in2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 500.110 596.000 500.390 600.000 ;
    END
  END in2[16]
  PIN in2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 506.090 596.000 506.370 600.000 ;
    END
  END in2[17]
  PIN in2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 512.070 596.000 512.350 600.000 ;
    END
  END in2[18]
  PIN in2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 518.050 596.000 518.330 600.000 ;
    END
  END in2[19]
  PIN in2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 410.410 596.000 410.690 600.000 ;
    END
  END in2[1]
  PIN in2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 524.030 596.000 524.310 600.000 ;
    END
  END in2[20]
  PIN in2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 530.010 596.000 530.290 600.000 ;
    END
  END in2[21]
  PIN in2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 535.990 596.000 536.270 600.000 ;
    END
  END in2[22]
  PIN in2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 541.970 596.000 542.250 600.000 ;
    END
  END in2[23]
  PIN in2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 547.950 596.000 548.230 600.000 ;
    END
  END in2[24]
  PIN in2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 553.930 596.000 554.210 600.000 ;
    END
  END in2[25]
  PIN in2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 596.000 560.190 600.000 ;
    END
  END in2[26]
  PIN in2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 565.890 596.000 566.170 600.000 ;
    END
  END in2[27]
  PIN in2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 571.870 596.000 572.150 600.000 ;
    END
  END in2[28]
  PIN in2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 577.850 596.000 578.130 600.000 ;
    END
  END in2[29]
  PIN in2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 416.390 596.000 416.670 600.000 ;
    END
  END in2[2]
  PIN in2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 583.830 596.000 584.110 600.000 ;
    END
  END in2[30]
  PIN in2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 589.810 596.000 590.090 600.000 ;
    END
  END in2[31]
  PIN in2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 422.370 596.000 422.650 600.000 ;
    END
  END in2[3]
  PIN in2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 596.000 428.630 600.000 ;
    END
  END in2[4]
  PIN in2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 434.330 596.000 434.610 600.000 ;
    END
  END in2[5]
  PIN in2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 440.310 596.000 440.590 600.000 ;
    END
  END in2[6]
  PIN in2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 446.290 596.000 446.570 600.000 ;
    END
  END in2[7]
  PIN in2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 452.270 596.000 452.550 600.000 ;
    END
  END in2[8]
  PIN in2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 458.250 596.000 458.530 600.000 ;
    END
  END in2[9]
  PIN out0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 40.840 600.000 41.440 ;
    END
  END out0[0]
  PIN out0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 95.240 600.000 95.840 ;
    END
  END out0[10]
  PIN out0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 100.680 600.000 101.280 ;
    END
  END out0[11]
  PIN out0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 106.120 600.000 106.720 ;
    END
  END out0[12]
  PIN out0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 111.560 600.000 112.160 ;
    END
  END out0[13]
  PIN out0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 117.000 600.000 117.600 ;
    END
  END out0[14]
  PIN out0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 122.440 600.000 123.040 ;
    END
  END out0[15]
  PIN out0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 127.880 600.000 128.480 ;
    END
  END out0[16]
  PIN out0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 133.320 600.000 133.920 ;
    END
  END out0[17]
  PIN out0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 138.760 600.000 139.360 ;
    END
  END out0[18]
  PIN out0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 144.200 600.000 144.800 ;
    END
  END out0[19]
  PIN out0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 46.280 600.000 46.880 ;
    END
  END out0[1]
  PIN out0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 149.640 600.000 150.240 ;
    END
  END out0[20]
  PIN out0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 155.080 600.000 155.680 ;
    END
  END out0[21]
  PIN out0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 160.520 600.000 161.120 ;
    END
  END out0[22]
  PIN out0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 165.960 600.000 166.560 ;
    END
  END out0[23]
  PIN out0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 171.400 600.000 172.000 ;
    END
  END out0[24]
  PIN out0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 176.840 600.000 177.440 ;
    END
  END out0[25]
  PIN out0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 182.280 600.000 182.880 ;
    END
  END out0[26]
  PIN out0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 187.720 600.000 188.320 ;
    END
  END out0[27]
  PIN out0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 193.160 600.000 193.760 ;
    END
  END out0[28]
  PIN out0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 198.600 600.000 199.200 ;
    END
  END out0[29]
  PIN out0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 51.720 600.000 52.320 ;
    END
  END out0[2]
  PIN out0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 204.040 600.000 204.640 ;
    END
  END out0[30]
  PIN out0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 209.480 600.000 210.080 ;
    END
  END out0[31]
  PIN out0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 57.160 600.000 57.760 ;
    END
  END out0[3]
  PIN out0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 62.600 600.000 63.200 ;
    END
  END out0[4]
  PIN out0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 68.040 600.000 68.640 ;
    END
  END out0[5]
  PIN out0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 73.480 600.000 74.080 ;
    END
  END out0[6]
  PIN out0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 78.920 600.000 79.520 ;
    END
  END out0[7]
  PIN out0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 84.360 600.000 84.960 ;
    END
  END out0[8]
  PIN out0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 89.800 600.000 90.400 ;
    END
  END out0[9]
  PIN out1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 214.920 600.000 215.520 ;
    END
  END out1[0]
  PIN out1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 269.320 600.000 269.920 ;
    END
  END out1[10]
  PIN out1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 274.760 600.000 275.360 ;
    END
  END out1[11]
  PIN out1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 280.200 600.000 280.800 ;
    END
  END out1[12]
  PIN out1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 285.640 600.000 286.240 ;
    END
  END out1[13]
  PIN out1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.080 600.000 291.680 ;
    END
  END out1[14]
  PIN out1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 296.520 600.000 297.120 ;
    END
  END out1[15]
  PIN out1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 301.960 600.000 302.560 ;
    END
  END out1[16]
  PIN out1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 307.400 600.000 308.000 ;
    END
  END out1[17]
  PIN out1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 312.840 600.000 313.440 ;
    END
  END out1[18]
  PIN out1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 318.280 600.000 318.880 ;
    END
  END out1[19]
  PIN out1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 220.360 600.000 220.960 ;
    END
  END out1[1]
  PIN out1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 323.720 600.000 324.320 ;
    END
  END out1[20]
  PIN out1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 329.160 600.000 329.760 ;
    END
  END out1[21]
  PIN out1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 334.600 600.000 335.200 ;
    END
  END out1[22]
  PIN out1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 340.040 600.000 340.640 ;
    END
  END out1[23]
  PIN out1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 345.480 600.000 346.080 ;
    END
  END out1[24]
  PIN out1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 350.920 600.000 351.520 ;
    END
  END out1[25]
  PIN out1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 356.360 600.000 356.960 ;
    END
  END out1[26]
  PIN out1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 361.800 600.000 362.400 ;
    END
  END out1[27]
  PIN out1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 367.240 600.000 367.840 ;
    END
  END out1[28]
  PIN out1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 372.680 600.000 373.280 ;
    END
  END out1[29]
  PIN out1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 225.800 600.000 226.400 ;
    END
  END out1[2]
  PIN out1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 378.120 600.000 378.720 ;
    END
  END out1[30]
  PIN out1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 383.560 600.000 384.160 ;
    END
  END out1[31]
  PIN out1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 231.240 600.000 231.840 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 236.680 600.000 237.280 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 242.120 600.000 242.720 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 247.560 600.000 248.160 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 253.000 600.000 253.600 ;
    END
  END out1[7]
  PIN out1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 258.440 600.000 259.040 ;
    END
  END out1[8]
  PIN out1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 263.880 600.000 264.480 ;
    END
  END out1[9]
  PIN out2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 389.000 600.000 389.600 ;
    END
  END out2[0]
  PIN out2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 443.400 600.000 444.000 ;
    END
  END out2[10]
  PIN out2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 448.840 600.000 449.440 ;
    END
  END out2[11]
  PIN out2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 454.280 600.000 454.880 ;
    END
  END out2[12]
  PIN out2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 459.720 600.000 460.320 ;
    END
  END out2[13]
  PIN out2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 465.160 600.000 465.760 ;
    END
  END out2[14]
  PIN out2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 470.600 600.000 471.200 ;
    END
  END out2[15]
  PIN out2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 476.040 600.000 476.640 ;
    END
  END out2[16]
  PIN out2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 481.480 600.000 482.080 ;
    END
  END out2[17]
  PIN out2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 486.920 600.000 487.520 ;
    END
  END out2[18]
  PIN out2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 492.360 600.000 492.960 ;
    END
  END out2[19]
  PIN out2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 394.440 600.000 395.040 ;
    END
  END out2[1]
  PIN out2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 497.800 600.000 498.400 ;
    END
  END out2[20]
  PIN out2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 503.240 600.000 503.840 ;
    END
  END out2[21]
  PIN out2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 508.680 600.000 509.280 ;
    END
  END out2[22]
  PIN out2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 514.120 600.000 514.720 ;
    END
  END out2[23]
  PIN out2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 519.560 600.000 520.160 ;
    END
  END out2[24]
  PIN out2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 525.000 600.000 525.600 ;
    END
  END out2[25]
  PIN out2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 530.440 600.000 531.040 ;
    END
  END out2[26]
  PIN out2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 535.880 600.000 536.480 ;
    END
  END out2[27]
  PIN out2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 541.320 600.000 541.920 ;
    END
  END out2[28]
  PIN out2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 546.760 600.000 547.360 ;
    END
  END out2[29]
  PIN out2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 399.880 600.000 400.480 ;
    END
  END out2[2]
  PIN out2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 552.200 600.000 552.800 ;
    END
  END out2[30]
  PIN out2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 557.640 600.000 558.240 ;
    END
  END out2[31]
  PIN out2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 405.320 600.000 405.920 ;
    END
  END out2[3]
  PIN out2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 410.760 600.000 411.360 ;
    END
  END out2[4]
  PIN out2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 416.200 600.000 416.800 ;
    END
  END out2[5]
  PIN out2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 421.640 600.000 422.240 ;
    END
  END out2[6]
  PIN out2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 427.080 600.000 427.680 ;
    END
  END out2[7]
  PIN out2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 432.520 600.000 433.120 ;
    END
  END out2[8]
  PIN out2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 437.960 600.000 438.560 ;
    END
  END out2[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 15.730 596.000 16.010 600.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 587.605 ;
      LAYER met1 ;
        RECT 1.450 0.720 598.390 595.640 ;
      LAYER met2 ;
        RECT 1.470 595.720 9.470 596.770 ;
        RECT 10.310 595.720 15.450 596.770 ;
        RECT 16.290 595.720 21.430 596.770 ;
        RECT 22.270 595.720 27.410 596.770 ;
        RECT 28.250 595.720 33.390 596.770 ;
        RECT 34.230 595.720 39.370 596.770 ;
        RECT 40.210 595.720 45.350 596.770 ;
        RECT 46.190 595.720 51.330 596.770 ;
        RECT 52.170 595.720 57.310 596.770 ;
        RECT 58.150 595.720 63.290 596.770 ;
        RECT 64.130 595.720 69.270 596.770 ;
        RECT 70.110 595.720 75.250 596.770 ;
        RECT 76.090 595.720 81.230 596.770 ;
        RECT 82.070 595.720 87.210 596.770 ;
        RECT 88.050 595.720 93.190 596.770 ;
        RECT 94.030 595.720 99.170 596.770 ;
        RECT 100.010 595.720 105.150 596.770 ;
        RECT 105.990 595.720 111.130 596.770 ;
        RECT 111.970 595.720 117.110 596.770 ;
        RECT 117.950 595.720 123.090 596.770 ;
        RECT 123.930 595.720 129.070 596.770 ;
        RECT 129.910 595.720 135.050 596.770 ;
        RECT 135.890 595.720 141.030 596.770 ;
        RECT 141.870 595.720 147.010 596.770 ;
        RECT 147.850 595.720 152.990 596.770 ;
        RECT 153.830 595.720 158.970 596.770 ;
        RECT 159.810 595.720 164.950 596.770 ;
        RECT 165.790 595.720 170.930 596.770 ;
        RECT 171.770 595.720 176.910 596.770 ;
        RECT 177.750 595.720 182.890 596.770 ;
        RECT 183.730 595.720 188.870 596.770 ;
        RECT 189.710 595.720 194.850 596.770 ;
        RECT 195.690 595.720 200.830 596.770 ;
        RECT 201.670 595.720 206.810 596.770 ;
        RECT 207.650 595.720 212.790 596.770 ;
        RECT 213.630 595.720 218.770 596.770 ;
        RECT 219.610 595.720 224.750 596.770 ;
        RECT 225.590 595.720 230.730 596.770 ;
        RECT 231.570 595.720 236.710 596.770 ;
        RECT 237.550 595.720 242.690 596.770 ;
        RECT 243.530 595.720 248.670 596.770 ;
        RECT 249.510 595.720 254.650 596.770 ;
        RECT 255.490 595.720 260.630 596.770 ;
        RECT 261.470 595.720 266.610 596.770 ;
        RECT 267.450 595.720 272.590 596.770 ;
        RECT 273.430 595.720 278.570 596.770 ;
        RECT 279.410 595.720 284.550 596.770 ;
        RECT 285.390 595.720 290.530 596.770 ;
        RECT 291.370 595.720 296.510 596.770 ;
        RECT 297.350 595.720 302.490 596.770 ;
        RECT 303.330 595.720 308.470 596.770 ;
        RECT 309.310 595.720 314.450 596.770 ;
        RECT 315.290 595.720 320.430 596.770 ;
        RECT 321.270 595.720 326.410 596.770 ;
        RECT 327.250 595.720 332.390 596.770 ;
        RECT 333.230 595.720 338.370 596.770 ;
        RECT 339.210 595.720 344.350 596.770 ;
        RECT 345.190 595.720 350.330 596.770 ;
        RECT 351.170 595.720 356.310 596.770 ;
        RECT 357.150 595.720 362.290 596.770 ;
        RECT 363.130 595.720 368.270 596.770 ;
        RECT 369.110 595.720 374.250 596.770 ;
        RECT 375.090 595.720 380.230 596.770 ;
        RECT 381.070 595.720 386.210 596.770 ;
        RECT 387.050 595.720 392.190 596.770 ;
        RECT 393.030 595.720 398.170 596.770 ;
        RECT 399.010 595.720 404.150 596.770 ;
        RECT 404.990 595.720 410.130 596.770 ;
        RECT 410.970 595.720 416.110 596.770 ;
        RECT 416.950 595.720 422.090 596.770 ;
        RECT 422.930 595.720 428.070 596.770 ;
        RECT 428.910 595.720 434.050 596.770 ;
        RECT 434.890 595.720 440.030 596.770 ;
        RECT 440.870 595.720 446.010 596.770 ;
        RECT 446.850 595.720 451.990 596.770 ;
        RECT 452.830 595.720 457.970 596.770 ;
        RECT 458.810 595.720 463.950 596.770 ;
        RECT 464.790 595.720 469.930 596.770 ;
        RECT 470.770 595.720 475.910 596.770 ;
        RECT 476.750 595.720 481.890 596.770 ;
        RECT 482.730 595.720 487.870 596.770 ;
        RECT 488.710 595.720 493.850 596.770 ;
        RECT 494.690 595.720 499.830 596.770 ;
        RECT 500.670 595.720 505.810 596.770 ;
        RECT 506.650 595.720 511.790 596.770 ;
        RECT 512.630 595.720 517.770 596.770 ;
        RECT 518.610 595.720 523.750 596.770 ;
        RECT 524.590 595.720 529.730 596.770 ;
        RECT 530.570 595.720 535.710 596.770 ;
        RECT 536.550 595.720 541.690 596.770 ;
        RECT 542.530 595.720 547.670 596.770 ;
        RECT 548.510 595.720 553.650 596.770 ;
        RECT 554.490 595.720 559.630 596.770 ;
        RECT 560.470 595.720 565.610 596.770 ;
        RECT 566.450 595.720 571.590 596.770 ;
        RECT 572.430 595.720 577.570 596.770 ;
        RECT 578.410 595.720 583.550 596.770 ;
        RECT 584.390 595.720 589.530 596.770 ;
        RECT 590.370 595.720 598.370 596.770 ;
        RECT 1.470 4.280 598.370 595.720 ;
        RECT 1.470 0.690 9.470 4.280 ;
        RECT 10.310 0.690 15.450 4.280 ;
        RECT 16.290 0.690 21.430 4.280 ;
        RECT 22.270 0.690 27.410 4.280 ;
        RECT 28.250 0.690 33.390 4.280 ;
        RECT 34.230 0.690 39.370 4.280 ;
        RECT 40.210 0.690 45.350 4.280 ;
        RECT 46.190 0.690 51.330 4.280 ;
        RECT 52.170 0.690 57.310 4.280 ;
        RECT 58.150 0.690 63.290 4.280 ;
        RECT 64.130 0.690 69.270 4.280 ;
        RECT 70.110 0.690 75.250 4.280 ;
        RECT 76.090 0.690 81.230 4.280 ;
        RECT 82.070 0.690 87.210 4.280 ;
        RECT 88.050 0.690 93.190 4.280 ;
        RECT 94.030 0.690 99.170 4.280 ;
        RECT 100.010 0.690 105.150 4.280 ;
        RECT 105.990 0.690 111.130 4.280 ;
        RECT 111.970 0.690 117.110 4.280 ;
        RECT 117.950 0.690 123.090 4.280 ;
        RECT 123.930 0.690 129.070 4.280 ;
        RECT 129.910 0.690 135.050 4.280 ;
        RECT 135.890 0.690 141.030 4.280 ;
        RECT 141.870 0.690 147.010 4.280 ;
        RECT 147.850 0.690 152.990 4.280 ;
        RECT 153.830 0.690 158.970 4.280 ;
        RECT 159.810 0.690 164.950 4.280 ;
        RECT 165.790 0.690 170.930 4.280 ;
        RECT 171.770 0.690 176.910 4.280 ;
        RECT 177.750 0.690 182.890 4.280 ;
        RECT 183.730 0.690 188.870 4.280 ;
        RECT 189.710 0.690 194.850 4.280 ;
        RECT 195.690 0.690 200.830 4.280 ;
        RECT 201.670 0.690 206.810 4.280 ;
        RECT 207.650 0.690 212.790 4.280 ;
        RECT 213.630 0.690 218.770 4.280 ;
        RECT 219.610 0.690 224.750 4.280 ;
        RECT 225.590 0.690 230.730 4.280 ;
        RECT 231.570 0.690 236.710 4.280 ;
        RECT 237.550 0.690 242.690 4.280 ;
        RECT 243.530 0.690 248.670 4.280 ;
        RECT 249.510 0.690 254.650 4.280 ;
        RECT 255.490 0.690 260.630 4.280 ;
        RECT 261.470 0.690 266.610 4.280 ;
        RECT 267.450 0.690 272.590 4.280 ;
        RECT 273.430 0.690 278.570 4.280 ;
        RECT 279.410 0.690 284.550 4.280 ;
        RECT 285.390 0.690 290.530 4.280 ;
        RECT 291.370 0.690 296.510 4.280 ;
        RECT 297.350 0.690 302.490 4.280 ;
        RECT 303.330 0.690 308.470 4.280 ;
        RECT 309.310 0.690 314.450 4.280 ;
        RECT 315.290 0.690 320.430 4.280 ;
        RECT 321.270 0.690 326.410 4.280 ;
        RECT 327.250 0.690 332.390 4.280 ;
        RECT 333.230 0.690 338.370 4.280 ;
        RECT 339.210 0.690 344.350 4.280 ;
        RECT 345.190 0.690 350.330 4.280 ;
        RECT 351.170 0.690 356.310 4.280 ;
        RECT 357.150 0.690 362.290 4.280 ;
        RECT 363.130 0.690 368.270 4.280 ;
        RECT 369.110 0.690 374.250 4.280 ;
        RECT 375.090 0.690 380.230 4.280 ;
        RECT 381.070 0.690 386.210 4.280 ;
        RECT 387.050 0.690 392.190 4.280 ;
        RECT 393.030 0.690 398.170 4.280 ;
        RECT 399.010 0.690 404.150 4.280 ;
        RECT 404.990 0.690 410.130 4.280 ;
        RECT 410.970 0.690 416.110 4.280 ;
        RECT 416.950 0.690 422.090 4.280 ;
        RECT 422.930 0.690 428.070 4.280 ;
        RECT 428.910 0.690 434.050 4.280 ;
        RECT 434.890 0.690 440.030 4.280 ;
        RECT 440.870 0.690 446.010 4.280 ;
        RECT 446.850 0.690 451.990 4.280 ;
        RECT 452.830 0.690 457.970 4.280 ;
        RECT 458.810 0.690 463.950 4.280 ;
        RECT 464.790 0.690 469.930 4.280 ;
        RECT 470.770 0.690 475.910 4.280 ;
        RECT 476.750 0.690 481.890 4.280 ;
        RECT 482.730 0.690 487.870 4.280 ;
        RECT 488.710 0.690 493.850 4.280 ;
        RECT 494.690 0.690 499.830 4.280 ;
        RECT 500.670 0.690 505.810 4.280 ;
        RECT 506.650 0.690 511.790 4.280 ;
        RECT 512.630 0.690 517.770 4.280 ;
        RECT 518.610 0.690 523.750 4.280 ;
        RECT 524.590 0.690 529.730 4.280 ;
        RECT 530.570 0.690 535.710 4.280 ;
        RECT 536.550 0.690 541.690 4.280 ;
        RECT 542.530 0.690 547.670 4.280 ;
        RECT 548.510 0.690 553.650 4.280 ;
        RECT 554.490 0.690 559.630 4.280 ;
        RECT 560.470 0.690 565.610 4.280 ;
        RECT 566.450 0.690 571.590 4.280 ;
        RECT 572.430 0.690 577.570 4.280 ;
        RECT 578.410 0.690 583.550 4.280 ;
        RECT 584.390 0.690 589.530 4.280 ;
        RECT 590.370 0.690 598.370 4.280 ;
      LAYER met3 ;
        RECT 1.445 561.360 598.395 587.685 ;
        RECT 4.400 559.960 598.395 561.360 ;
        RECT 1.445 558.640 598.395 559.960 ;
        RECT 1.445 557.240 595.600 558.640 ;
        RECT 1.445 553.200 598.395 557.240 ;
        RECT 4.400 551.800 595.600 553.200 ;
        RECT 1.445 547.760 598.395 551.800 ;
        RECT 1.445 546.360 595.600 547.760 ;
        RECT 1.445 545.040 598.395 546.360 ;
        RECT 4.400 543.640 598.395 545.040 ;
        RECT 1.445 542.320 598.395 543.640 ;
        RECT 1.445 540.920 595.600 542.320 ;
        RECT 1.445 536.880 598.395 540.920 ;
        RECT 4.400 535.480 595.600 536.880 ;
        RECT 1.445 531.440 598.395 535.480 ;
        RECT 1.445 530.040 595.600 531.440 ;
        RECT 1.445 528.720 598.395 530.040 ;
        RECT 4.400 527.320 598.395 528.720 ;
        RECT 1.445 526.000 598.395 527.320 ;
        RECT 1.445 524.600 595.600 526.000 ;
        RECT 1.445 520.560 598.395 524.600 ;
        RECT 4.400 519.160 595.600 520.560 ;
        RECT 1.445 515.120 598.395 519.160 ;
        RECT 1.445 513.720 595.600 515.120 ;
        RECT 1.445 512.400 598.395 513.720 ;
        RECT 4.400 511.000 598.395 512.400 ;
        RECT 1.445 509.680 598.395 511.000 ;
        RECT 1.445 508.280 595.600 509.680 ;
        RECT 1.445 504.240 598.395 508.280 ;
        RECT 4.400 502.840 595.600 504.240 ;
        RECT 1.445 498.800 598.395 502.840 ;
        RECT 1.445 497.400 595.600 498.800 ;
        RECT 1.445 496.080 598.395 497.400 ;
        RECT 4.400 494.680 598.395 496.080 ;
        RECT 1.445 493.360 598.395 494.680 ;
        RECT 1.445 491.960 595.600 493.360 ;
        RECT 1.445 487.920 598.395 491.960 ;
        RECT 4.400 486.520 595.600 487.920 ;
        RECT 1.445 482.480 598.395 486.520 ;
        RECT 1.445 481.080 595.600 482.480 ;
        RECT 1.445 479.760 598.395 481.080 ;
        RECT 4.400 478.360 598.395 479.760 ;
        RECT 1.445 477.040 598.395 478.360 ;
        RECT 1.445 475.640 595.600 477.040 ;
        RECT 1.445 471.600 598.395 475.640 ;
        RECT 4.400 470.200 595.600 471.600 ;
        RECT 1.445 466.160 598.395 470.200 ;
        RECT 1.445 464.760 595.600 466.160 ;
        RECT 1.445 463.440 598.395 464.760 ;
        RECT 4.400 462.040 598.395 463.440 ;
        RECT 1.445 460.720 598.395 462.040 ;
        RECT 1.445 459.320 595.600 460.720 ;
        RECT 1.445 455.280 598.395 459.320 ;
        RECT 4.400 453.880 595.600 455.280 ;
        RECT 1.445 449.840 598.395 453.880 ;
        RECT 1.445 448.440 595.600 449.840 ;
        RECT 1.445 447.120 598.395 448.440 ;
        RECT 4.400 445.720 598.395 447.120 ;
        RECT 1.445 444.400 598.395 445.720 ;
        RECT 1.445 443.000 595.600 444.400 ;
        RECT 1.445 438.960 598.395 443.000 ;
        RECT 4.400 437.560 595.600 438.960 ;
        RECT 1.445 433.520 598.395 437.560 ;
        RECT 1.445 432.120 595.600 433.520 ;
        RECT 1.445 430.800 598.395 432.120 ;
        RECT 4.400 429.400 598.395 430.800 ;
        RECT 1.445 428.080 598.395 429.400 ;
        RECT 1.445 426.680 595.600 428.080 ;
        RECT 1.445 422.640 598.395 426.680 ;
        RECT 4.400 421.240 595.600 422.640 ;
        RECT 1.445 417.200 598.395 421.240 ;
        RECT 1.445 415.800 595.600 417.200 ;
        RECT 1.445 414.480 598.395 415.800 ;
        RECT 4.400 413.080 598.395 414.480 ;
        RECT 1.445 411.760 598.395 413.080 ;
        RECT 1.445 410.360 595.600 411.760 ;
        RECT 1.445 406.320 598.395 410.360 ;
        RECT 4.400 404.920 595.600 406.320 ;
        RECT 1.445 400.880 598.395 404.920 ;
        RECT 1.445 399.480 595.600 400.880 ;
        RECT 1.445 398.160 598.395 399.480 ;
        RECT 4.400 396.760 598.395 398.160 ;
        RECT 1.445 395.440 598.395 396.760 ;
        RECT 1.445 394.040 595.600 395.440 ;
        RECT 1.445 390.000 598.395 394.040 ;
        RECT 4.400 388.600 595.600 390.000 ;
        RECT 1.445 384.560 598.395 388.600 ;
        RECT 1.445 383.160 595.600 384.560 ;
        RECT 1.445 381.840 598.395 383.160 ;
        RECT 4.400 380.440 598.395 381.840 ;
        RECT 1.445 379.120 598.395 380.440 ;
        RECT 1.445 377.720 595.600 379.120 ;
        RECT 1.445 373.680 598.395 377.720 ;
        RECT 4.400 372.280 595.600 373.680 ;
        RECT 1.445 368.240 598.395 372.280 ;
        RECT 1.445 366.840 595.600 368.240 ;
        RECT 1.445 365.520 598.395 366.840 ;
        RECT 4.400 364.120 598.395 365.520 ;
        RECT 1.445 362.800 598.395 364.120 ;
        RECT 1.445 361.400 595.600 362.800 ;
        RECT 1.445 357.360 598.395 361.400 ;
        RECT 4.400 355.960 595.600 357.360 ;
        RECT 1.445 351.920 598.395 355.960 ;
        RECT 1.445 350.520 595.600 351.920 ;
        RECT 1.445 349.200 598.395 350.520 ;
        RECT 4.400 347.800 598.395 349.200 ;
        RECT 1.445 346.480 598.395 347.800 ;
        RECT 1.445 345.080 595.600 346.480 ;
        RECT 1.445 341.040 598.395 345.080 ;
        RECT 4.400 339.640 595.600 341.040 ;
        RECT 1.445 335.600 598.395 339.640 ;
        RECT 1.445 334.200 595.600 335.600 ;
        RECT 1.445 332.880 598.395 334.200 ;
        RECT 4.400 331.480 598.395 332.880 ;
        RECT 1.445 330.160 598.395 331.480 ;
        RECT 1.445 328.760 595.600 330.160 ;
        RECT 1.445 324.720 598.395 328.760 ;
        RECT 4.400 323.320 595.600 324.720 ;
        RECT 1.445 319.280 598.395 323.320 ;
        RECT 1.445 317.880 595.600 319.280 ;
        RECT 1.445 316.560 598.395 317.880 ;
        RECT 4.400 315.160 598.395 316.560 ;
        RECT 1.445 313.840 598.395 315.160 ;
        RECT 1.445 312.440 595.600 313.840 ;
        RECT 1.445 308.400 598.395 312.440 ;
        RECT 4.400 307.000 595.600 308.400 ;
        RECT 1.445 302.960 598.395 307.000 ;
        RECT 1.445 301.560 595.600 302.960 ;
        RECT 1.445 300.240 598.395 301.560 ;
        RECT 4.400 298.840 598.395 300.240 ;
        RECT 1.445 297.520 598.395 298.840 ;
        RECT 1.445 296.120 595.600 297.520 ;
        RECT 1.445 292.080 598.395 296.120 ;
        RECT 4.400 290.680 595.600 292.080 ;
        RECT 1.445 286.640 598.395 290.680 ;
        RECT 1.445 285.240 595.600 286.640 ;
        RECT 1.445 283.920 598.395 285.240 ;
        RECT 4.400 282.520 598.395 283.920 ;
        RECT 1.445 281.200 598.395 282.520 ;
        RECT 1.445 279.800 595.600 281.200 ;
        RECT 1.445 275.760 598.395 279.800 ;
        RECT 4.400 274.360 595.600 275.760 ;
        RECT 1.445 270.320 598.395 274.360 ;
        RECT 1.445 268.920 595.600 270.320 ;
        RECT 1.445 267.600 598.395 268.920 ;
        RECT 4.400 266.200 598.395 267.600 ;
        RECT 1.445 264.880 598.395 266.200 ;
        RECT 1.445 263.480 595.600 264.880 ;
        RECT 1.445 259.440 598.395 263.480 ;
        RECT 4.400 258.040 595.600 259.440 ;
        RECT 1.445 254.000 598.395 258.040 ;
        RECT 1.445 252.600 595.600 254.000 ;
        RECT 1.445 251.280 598.395 252.600 ;
        RECT 4.400 249.880 598.395 251.280 ;
        RECT 1.445 248.560 598.395 249.880 ;
        RECT 1.445 247.160 595.600 248.560 ;
        RECT 1.445 243.120 598.395 247.160 ;
        RECT 4.400 241.720 595.600 243.120 ;
        RECT 1.445 237.680 598.395 241.720 ;
        RECT 1.445 236.280 595.600 237.680 ;
        RECT 1.445 234.960 598.395 236.280 ;
        RECT 4.400 233.560 598.395 234.960 ;
        RECT 1.445 232.240 598.395 233.560 ;
        RECT 1.445 230.840 595.600 232.240 ;
        RECT 1.445 226.800 598.395 230.840 ;
        RECT 4.400 225.400 595.600 226.800 ;
        RECT 1.445 221.360 598.395 225.400 ;
        RECT 1.445 219.960 595.600 221.360 ;
        RECT 1.445 218.640 598.395 219.960 ;
        RECT 4.400 217.240 598.395 218.640 ;
        RECT 1.445 215.920 598.395 217.240 ;
        RECT 1.445 214.520 595.600 215.920 ;
        RECT 1.445 210.480 598.395 214.520 ;
        RECT 4.400 209.080 595.600 210.480 ;
        RECT 1.445 205.040 598.395 209.080 ;
        RECT 1.445 203.640 595.600 205.040 ;
        RECT 1.445 202.320 598.395 203.640 ;
        RECT 4.400 200.920 598.395 202.320 ;
        RECT 1.445 199.600 598.395 200.920 ;
        RECT 1.445 198.200 595.600 199.600 ;
        RECT 1.445 194.160 598.395 198.200 ;
        RECT 4.400 192.760 595.600 194.160 ;
        RECT 1.445 188.720 598.395 192.760 ;
        RECT 1.445 187.320 595.600 188.720 ;
        RECT 1.445 186.000 598.395 187.320 ;
        RECT 4.400 184.600 598.395 186.000 ;
        RECT 1.445 183.280 598.395 184.600 ;
        RECT 1.445 181.880 595.600 183.280 ;
        RECT 1.445 177.840 598.395 181.880 ;
        RECT 4.400 176.440 595.600 177.840 ;
        RECT 1.445 172.400 598.395 176.440 ;
        RECT 1.445 171.000 595.600 172.400 ;
        RECT 1.445 169.680 598.395 171.000 ;
        RECT 4.400 168.280 598.395 169.680 ;
        RECT 1.445 166.960 598.395 168.280 ;
        RECT 1.445 165.560 595.600 166.960 ;
        RECT 1.445 161.520 598.395 165.560 ;
        RECT 4.400 160.120 595.600 161.520 ;
        RECT 1.445 156.080 598.395 160.120 ;
        RECT 1.445 154.680 595.600 156.080 ;
        RECT 1.445 153.360 598.395 154.680 ;
        RECT 4.400 151.960 598.395 153.360 ;
        RECT 1.445 150.640 598.395 151.960 ;
        RECT 1.445 149.240 595.600 150.640 ;
        RECT 1.445 145.200 598.395 149.240 ;
        RECT 4.400 143.800 595.600 145.200 ;
        RECT 1.445 139.760 598.395 143.800 ;
        RECT 1.445 138.360 595.600 139.760 ;
        RECT 1.445 137.040 598.395 138.360 ;
        RECT 4.400 135.640 598.395 137.040 ;
        RECT 1.445 134.320 598.395 135.640 ;
        RECT 1.445 132.920 595.600 134.320 ;
        RECT 1.445 128.880 598.395 132.920 ;
        RECT 4.400 127.480 595.600 128.880 ;
        RECT 1.445 123.440 598.395 127.480 ;
        RECT 1.445 122.040 595.600 123.440 ;
        RECT 1.445 120.720 598.395 122.040 ;
        RECT 4.400 119.320 598.395 120.720 ;
        RECT 1.445 118.000 598.395 119.320 ;
        RECT 1.445 116.600 595.600 118.000 ;
        RECT 1.445 112.560 598.395 116.600 ;
        RECT 4.400 111.160 595.600 112.560 ;
        RECT 1.445 107.120 598.395 111.160 ;
        RECT 1.445 105.720 595.600 107.120 ;
        RECT 1.445 104.400 598.395 105.720 ;
        RECT 4.400 103.000 598.395 104.400 ;
        RECT 1.445 101.680 598.395 103.000 ;
        RECT 1.445 100.280 595.600 101.680 ;
        RECT 1.445 96.240 598.395 100.280 ;
        RECT 4.400 94.840 595.600 96.240 ;
        RECT 1.445 90.800 598.395 94.840 ;
        RECT 1.445 89.400 595.600 90.800 ;
        RECT 1.445 88.080 598.395 89.400 ;
        RECT 4.400 86.680 598.395 88.080 ;
        RECT 1.445 85.360 598.395 86.680 ;
        RECT 1.445 83.960 595.600 85.360 ;
        RECT 1.445 79.920 598.395 83.960 ;
        RECT 4.400 78.520 595.600 79.920 ;
        RECT 1.445 74.480 598.395 78.520 ;
        RECT 1.445 73.080 595.600 74.480 ;
        RECT 1.445 71.760 598.395 73.080 ;
        RECT 4.400 70.360 598.395 71.760 ;
        RECT 1.445 69.040 598.395 70.360 ;
        RECT 1.445 67.640 595.600 69.040 ;
        RECT 1.445 63.600 598.395 67.640 ;
        RECT 4.400 62.200 595.600 63.600 ;
        RECT 1.445 58.160 598.395 62.200 ;
        RECT 1.445 56.760 595.600 58.160 ;
        RECT 1.445 55.440 598.395 56.760 ;
        RECT 4.400 54.040 598.395 55.440 ;
        RECT 1.445 52.720 598.395 54.040 ;
        RECT 1.445 51.320 595.600 52.720 ;
        RECT 1.445 47.280 598.395 51.320 ;
        RECT 4.400 45.880 595.600 47.280 ;
        RECT 1.445 41.840 598.395 45.880 ;
        RECT 1.445 40.440 595.600 41.840 ;
        RECT 1.445 39.120 598.395 40.440 ;
        RECT 4.400 37.720 598.395 39.120 ;
        RECT 1.445 2.895 598.395 37.720 ;
      LAYER met4 ;
        RECT 3.975 10.240 20.640 573.065 ;
        RECT 23.040 10.240 97.440 573.065 ;
        RECT 99.840 10.240 174.240 573.065 ;
        RECT 176.640 10.240 251.040 573.065 ;
        RECT 253.440 10.240 327.840 573.065 ;
        RECT 330.240 10.240 404.640 573.065 ;
        RECT 407.040 10.240 481.440 573.065 ;
        RECT 483.840 10.240 558.240 573.065 ;
        RECT 560.640 10.240 585.745 573.065 ;
        RECT 3.975 2.895 585.745 10.240 ;
  END
END Proc
END LIBRARY


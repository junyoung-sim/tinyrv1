`ifndef PROCDPATH_V
`define PROCDPATH_V

module ProcDpath
(
  
);



endmodule

`endif
magic
tech sky130A
magscale 1 2
timestamp 1740540685
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 290 144 119678 119128
<< metal2 >>
rect 1950 119200 2006 120000
rect 3146 119200 3202 120000
rect 4342 119200 4398 120000
rect 5538 119200 5594 120000
rect 6734 119200 6790 120000
rect 7930 119200 7986 120000
rect 9126 119200 9182 120000
rect 10322 119200 10378 120000
rect 11518 119200 11574 120000
rect 12714 119200 12770 120000
rect 13910 119200 13966 120000
rect 15106 119200 15162 120000
rect 16302 119200 16358 120000
rect 17498 119200 17554 120000
rect 18694 119200 18750 120000
rect 19890 119200 19946 120000
rect 21086 119200 21142 120000
rect 22282 119200 22338 120000
rect 23478 119200 23534 120000
rect 24674 119200 24730 120000
rect 25870 119200 25926 120000
rect 27066 119200 27122 120000
rect 28262 119200 28318 120000
rect 29458 119200 29514 120000
rect 30654 119200 30710 120000
rect 31850 119200 31906 120000
rect 33046 119200 33102 120000
rect 34242 119200 34298 120000
rect 35438 119200 35494 120000
rect 36634 119200 36690 120000
rect 37830 119200 37886 120000
rect 39026 119200 39082 120000
rect 40222 119200 40278 120000
rect 41418 119200 41474 120000
rect 42614 119200 42670 120000
rect 43810 119200 43866 120000
rect 45006 119200 45062 120000
rect 46202 119200 46258 120000
rect 47398 119200 47454 120000
rect 48594 119200 48650 120000
rect 49790 119200 49846 120000
rect 50986 119200 51042 120000
rect 52182 119200 52238 120000
rect 53378 119200 53434 120000
rect 54574 119200 54630 120000
rect 55770 119200 55826 120000
rect 56966 119200 57022 120000
rect 58162 119200 58218 120000
rect 59358 119200 59414 120000
rect 60554 119200 60610 120000
rect 61750 119200 61806 120000
rect 62946 119200 63002 120000
rect 64142 119200 64198 120000
rect 65338 119200 65394 120000
rect 66534 119200 66590 120000
rect 67730 119200 67786 120000
rect 68926 119200 68982 120000
rect 70122 119200 70178 120000
rect 71318 119200 71374 120000
rect 72514 119200 72570 120000
rect 73710 119200 73766 120000
rect 74906 119200 74962 120000
rect 76102 119200 76158 120000
rect 77298 119200 77354 120000
rect 78494 119200 78550 120000
rect 79690 119200 79746 120000
rect 80886 119200 80942 120000
rect 82082 119200 82138 120000
rect 83278 119200 83334 120000
rect 84474 119200 84530 120000
rect 85670 119200 85726 120000
rect 86866 119200 86922 120000
rect 88062 119200 88118 120000
rect 89258 119200 89314 120000
rect 90454 119200 90510 120000
rect 91650 119200 91706 120000
rect 92846 119200 92902 120000
rect 94042 119200 94098 120000
rect 95238 119200 95294 120000
rect 96434 119200 96490 120000
rect 97630 119200 97686 120000
rect 98826 119200 98882 120000
rect 100022 119200 100078 120000
rect 101218 119200 101274 120000
rect 102414 119200 102470 120000
rect 103610 119200 103666 120000
rect 104806 119200 104862 120000
rect 106002 119200 106058 120000
rect 107198 119200 107254 120000
rect 108394 119200 108450 120000
rect 109590 119200 109646 120000
rect 110786 119200 110842 120000
rect 111982 119200 112038 120000
rect 113178 119200 113234 120000
rect 114374 119200 114430 120000
rect 115570 119200 115626 120000
rect 116766 119200 116822 120000
rect 117962 119200 118018 120000
rect 1950 0 2006 800
rect 3146 0 3202 800
rect 4342 0 4398 800
rect 5538 0 5594 800
rect 6734 0 6790 800
rect 7930 0 7986 800
rect 9126 0 9182 800
rect 10322 0 10378 800
rect 11518 0 11574 800
rect 12714 0 12770 800
rect 13910 0 13966 800
rect 15106 0 15162 800
rect 16302 0 16358 800
rect 17498 0 17554 800
rect 18694 0 18750 800
rect 19890 0 19946 800
rect 21086 0 21142 800
rect 22282 0 22338 800
rect 23478 0 23534 800
rect 24674 0 24730 800
rect 25870 0 25926 800
rect 27066 0 27122 800
rect 28262 0 28318 800
rect 29458 0 29514 800
rect 30654 0 30710 800
rect 31850 0 31906 800
rect 33046 0 33102 800
rect 34242 0 34298 800
rect 35438 0 35494 800
rect 36634 0 36690 800
rect 37830 0 37886 800
rect 39026 0 39082 800
rect 40222 0 40278 800
rect 41418 0 41474 800
rect 42614 0 42670 800
rect 43810 0 43866 800
rect 45006 0 45062 800
rect 46202 0 46258 800
rect 47398 0 47454 800
rect 48594 0 48650 800
rect 49790 0 49846 800
rect 50986 0 51042 800
rect 52182 0 52238 800
rect 53378 0 53434 800
rect 54574 0 54630 800
rect 55770 0 55826 800
rect 56966 0 57022 800
rect 58162 0 58218 800
rect 59358 0 59414 800
rect 60554 0 60610 800
rect 61750 0 61806 800
rect 62946 0 63002 800
rect 64142 0 64198 800
rect 65338 0 65394 800
rect 66534 0 66590 800
rect 67730 0 67786 800
rect 68926 0 68982 800
rect 70122 0 70178 800
rect 71318 0 71374 800
rect 72514 0 72570 800
rect 73710 0 73766 800
rect 74906 0 74962 800
rect 76102 0 76158 800
rect 77298 0 77354 800
rect 78494 0 78550 800
rect 79690 0 79746 800
rect 80886 0 80942 800
rect 82082 0 82138 800
rect 83278 0 83334 800
rect 84474 0 84530 800
rect 85670 0 85726 800
rect 86866 0 86922 800
rect 88062 0 88118 800
rect 89258 0 89314 800
rect 90454 0 90510 800
rect 91650 0 91706 800
rect 92846 0 92902 800
rect 94042 0 94098 800
rect 95238 0 95294 800
rect 96434 0 96490 800
rect 97630 0 97686 800
rect 98826 0 98882 800
rect 100022 0 100078 800
rect 101218 0 101274 800
rect 102414 0 102470 800
rect 103610 0 103666 800
rect 104806 0 104862 800
rect 106002 0 106058 800
rect 107198 0 107254 800
rect 108394 0 108450 800
rect 109590 0 109646 800
rect 110786 0 110842 800
rect 111982 0 112038 800
rect 113178 0 113234 800
rect 114374 0 114430 800
rect 115570 0 115626 800
rect 116766 0 116822 800
rect 117962 0 118018 800
<< obsm2 >>
rect 294 119144 1894 119354
rect 2062 119144 3090 119354
rect 3258 119144 4286 119354
rect 4454 119144 5482 119354
rect 5650 119144 6678 119354
rect 6846 119144 7874 119354
rect 8042 119144 9070 119354
rect 9238 119144 10266 119354
rect 10434 119144 11462 119354
rect 11630 119144 12658 119354
rect 12826 119144 13854 119354
rect 14022 119144 15050 119354
rect 15218 119144 16246 119354
rect 16414 119144 17442 119354
rect 17610 119144 18638 119354
rect 18806 119144 19834 119354
rect 20002 119144 21030 119354
rect 21198 119144 22226 119354
rect 22394 119144 23422 119354
rect 23590 119144 24618 119354
rect 24786 119144 25814 119354
rect 25982 119144 27010 119354
rect 27178 119144 28206 119354
rect 28374 119144 29402 119354
rect 29570 119144 30598 119354
rect 30766 119144 31794 119354
rect 31962 119144 32990 119354
rect 33158 119144 34186 119354
rect 34354 119144 35382 119354
rect 35550 119144 36578 119354
rect 36746 119144 37774 119354
rect 37942 119144 38970 119354
rect 39138 119144 40166 119354
rect 40334 119144 41362 119354
rect 41530 119144 42558 119354
rect 42726 119144 43754 119354
rect 43922 119144 44950 119354
rect 45118 119144 46146 119354
rect 46314 119144 47342 119354
rect 47510 119144 48538 119354
rect 48706 119144 49734 119354
rect 49902 119144 50930 119354
rect 51098 119144 52126 119354
rect 52294 119144 53322 119354
rect 53490 119144 54518 119354
rect 54686 119144 55714 119354
rect 55882 119144 56910 119354
rect 57078 119144 58106 119354
rect 58274 119144 59302 119354
rect 59470 119144 60498 119354
rect 60666 119144 61694 119354
rect 61862 119144 62890 119354
rect 63058 119144 64086 119354
rect 64254 119144 65282 119354
rect 65450 119144 66478 119354
rect 66646 119144 67674 119354
rect 67842 119144 68870 119354
rect 69038 119144 70066 119354
rect 70234 119144 71262 119354
rect 71430 119144 72458 119354
rect 72626 119144 73654 119354
rect 73822 119144 74850 119354
rect 75018 119144 76046 119354
rect 76214 119144 77242 119354
rect 77410 119144 78438 119354
rect 78606 119144 79634 119354
rect 79802 119144 80830 119354
rect 80998 119144 82026 119354
rect 82194 119144 83222 119354
rect 83390 119144 84418 119354
rect 84586 119144 85614 119354
rect 85782 119144 86810 119354
rect 86978 119144 88006 119354
rect 88174 119144 89202 119354
rect 89370 119144 90398 119354
rect 90566 119144 91594 119354
rect 91762 119144 92790 119354
rect 92958 119144 93986 119354
rect 94154 119144 95182 119354
rect 95350 119144 96378 119354
rect 96546 119144 97574 119354
rect 97742 119144 98770 119354
rect 98938 119144 99966 119354
rect 100134 119144 101162 119354
rect 101330 119144 102358 119354
rect 102526 119144 103554 119354
rect 103722 119144 104750 119354
rect 104918 119144 105946 119354
rect 106114 119144 107142 119354
rect 107310 119144 108338 119354
rect 108506 119144 109534 119354
rect 109702 119144 110730 119354
rect 110898 119144 111926 119354
rect 112094 119144 113122 119354
rect 113290 119144 114318 119354
rect 114486 119144 115514 119354
rect 115682 119144 116710 119354
rect 116878 119144 117906 119354
rect 118074 119144 119674 119354
rect 294 856 119674 119144
rect 294 138 1894 856
rect 2062 138 3090 856
rect 3258 138 4286 856
rect 4454 138 5482 856
rect 5650 138 6678 856
rect 6846 138 7874 856
rect 8042 138 9070 856
rect 9238 138 10266 856
rect 10434 138 11462 856
rect 11630 138 12658 856
rect 12826 138 13854 856
rect 14022 138 15050 856
rect 15218 138 16246 856
rect 16414 138 17442 856
rect 17610 138 18638 856
rect 18806 138 19834 856
rect 20002 138 21030 856
rect 21198 138 22226 856
rect 22394 138 23422 856
rect 23590 138 24618 856
rect 24786 138 25814 856
rect 25982 138 27010 856
rect 27178 138 28206 856
rect 28374 138 29402 856
rect 29570 138 30598 856
rect 30766 138 31794 856
rect 31962 138 32990 856
rect 33158 138 34186 856
rect 34354 138 35382 856
rect 35550 138 36578 856
rect 36746 138 37774 856
rect 37942 138 38970 856
rect 39138 138 40166 856
rect 40334 138 41362 856
rect 41530 138 42558 856
rect 42726 138 43754 856
rect 43922 138 44950 856
rect 45118 138 46146 856
rect 46314 138 47342 856
rect 47510 138 48538 856
rect 48706 138 49734 856
rect 49902 138 50930 856
rect 51098 138 52126 856
rect 52294 138 53322 856
rect 53490 138 54518 856
rect 54686 138 55714 856
rect 55882 138 56910 856
rect 57078 138 58106 856
rect 58274 138 59302 856
rect 59470 138 60498 856
rect 60666 138 61694 856
rect 61862 138 62890 856
rect 63058 138 64086 856
rect 64254 138 65282 856
rect 65450 138 66478 856
rect 66646 138 67674 856
rect 67842 138 68870 856
rect 69038 138 70066 856
rect 70234 138 71262 856
rect 71430 138 72458 856
rect 72626 138 73654 856
rect 73822 138 74850 856
rect 75018 138 76046 856
rect 76214 138 77242 856
rect 77410 138 78438 856
rect 78606 138 79634 856
rect 79802 138 80830 856
rect 80998 138 82026 856
rect 82194 138 83222 856
rect 83390 138 84418 856
rect 84586 138 85614 856
rect 85782 138 86810 856
rect 86978 138 88006 856
rect 88174 138 89202 856
rect 89370 138 90398 856
rect 90566 138 91594 856
rect 91762 138 92790 856
rect 92958 138 93986 856
rect 94154 138 95182 856
rect 95350 138 96378 856
rect 96546 138 97574 856
rect 97742 138 98770 856
rect 98938 138 99966 856
rect 100134 138 101162 856
rect 101330 138 102358 856
rect 102526 138 103554 856
rect 103722 138 104750 856
rect 104918 138 105946 856
rect 106114 138 107142 856
rect 107310 138 108338 856
rect 108506 138 109534 856
rect 109702 138 110730 856
rect 110898 138 111926 856
rect 112094 138 113122 856
rect 113290 138 114318 856
rect 114486 138 115514 856
rect 115682 138 116710 856
rect 116878 138 117906 856
rect 118074 138 119674 856
<< metal3 >>
rect 0 112072 800 112192
rect 119200 111528 120000 111648
rect 0 110440 800 110560
rect 119200 110440 120000 110560
rect 119200 109352 120000 109472
rect 0 108808 800 108928
rect 119200 108264 120000 108384
rect 0 107176 800 107296
rect 119200 107176 120000 107296
rect 119200 106088 120000 106208
rect 0 105544 800 105664
rect 119200 105000 120000 105120
rect 0 103912 800 104032
rect 119200 103912 120000 104032
rect 119200 102824 120000 102944
rect 0 102280 800 102400
rect 119200 101736 120000 101856
rect 0 100648 800 100768
rect 119200 100648 120000 100768
rect 119200 99560 120000 99680
rect 0 99016 800 99136
rect 119200 98472 120000 98592
rect 0 97384 800 97504
rect 119200 97384 120000 97504
rect 119200 96296 120000 96416
rect 0 95752 800 95872
rect 119200 95208 120000 95328
rect 0 94120 800 94240
rect 119200 94120 120000 94240
rect 119200 93032 120000 93152
rect 0 92488 800 92608
rect 119200 91944 120000 92064
rect 0 90856 800 90976
rect 119200 90856 120000 90976
rect 119200 89768 120000 89888
rect 0 89224 800 89344
rect 119200 88680 120000 88800
rect 0 87592 800 87712
rect 119200 87592 120000 87712
rect 119200 86504 120000 86624
rect 0 85960 800 86080
rect 119200 85416 120000 85536
rect 0 84328 800 84448
rect 119200 84328 120000 84448
rect 119200 83240 120000 83360
rect 0 82696 800 82816
rect 119200 82152 120000 82272
rect 0 81064 800 81184
rect 119200 81064 120000 81184
rect 119200 79976 120000 80096
rect 0 79432 800 79552
rect 119200 78888 120000 79008
rect 0 77800 800 77920
rect 119200 77800 120000 77920
rect 119200 76712 120000 76832
rect 0 76168 800 76288
rect 119200 75624 120000 75744
rect 0 74536 800 74656
rect 119200 74536 120000 74656
rect 119200 73448 120000 73568
rect 0 72904 800 73024
rect 119200 72360 120000 72480
rect 0 71272 800 71392
rect 119200 71272 120000 71392
rect 119200 70184 120000 70304
rect 0 69640 800 69760
rect 119200 69096 120000 69216
rect 0 68008 800 68128
rect 119200 68008 120000 68128
rect 119200 66920 120000 67040
rect 0 66376 800 66496
rect 119200 65832 120000 65952
rect 0 64744 800 64864
rect 119200 64744 120000 64864
rect 119200 63656 120000 63776
rect 0 63112 800 63232
rect 119200 62568 120000 62688
rect 0 61480 800 61600
rect 119200 61480 120000 61600
rect 119200 60392 120000 60512
rect 0 59848 800 59968
rect 119200 59304 120000 59424
rect 0 58216 800 58336
rect 119200 58216 120000 58336
rect 119200 57128 120000 57248
rect 0 56584 800 56704
rect 119200 56040 120000 56160
rect 0 54952 800 55072
rect 119200 54952 120000 55072
rect 119200 53864 120000 53984
rect 0 53320 800 53440
rect 119200 52776 120000 52896
rect 0 51688 800 51808
rect 119200 51688 120000 51808
rect 119200 50600 120000 50720
rect 0 50056 800 50176
rect 119200 49512 120000 49632
rect 0 48424 800 48544
rect 119200 48424 120000 48544
rect 119200 47336 120000 47456
rect 0 46792 800 46912
rect 119200 46248 120000 46368
rect 0 45160 800 45280
rect 119200 45160 120000 45280
rect 119200 44072 120000 44192
rect 0 43528 800 43648
rect 119200 42984 120000 43104
rect 0 41896 800 42016
rect 119200 41896 120000 42016
rect 119200 40808 120000 40928
rect 0 40264 800 40384
rect 119200 39720 120000 39840
rect 0 38632 800 38752
rect 119200 38632 120000 38752
rect 119200 37544 120000 37664
rect 0 37000 800 37120
rect 119200 36456 120000 36576
rect 0 35368 800 35488
rect 119200 35368 120000 35488
rect 119200 34280 120000 34400
rect 0 33736 800 33856
rect 119200 33192 120000 33312
rect 0 32104 800 32224
rect 119200 32104 120000 32224
rect 119200 31016 120000 31136
rect 0 30472 800 30592
rect 119200 29928 120000 30048
rect 0 28840 800 28960
rect 119200 28840 120000 28960
rect 119200 27752 120000 27872
rect 0 27208 800 27328
rect 119200 26664 120000 26784
rect 0 25576 800 25696
rect 119200 25576 120000 25696
rect 119200 24488 120000 24608
rect 0 23944 800 24064
rect 119200 23400 120000 23520
rect 0 22312 800 22432
rect 119200 22312 120000 22432
rect 119200 21224 120000 21344
rect 0 20680 800 20800
rect 119200 20136 120000 20256
rect 0 19048 800 19168
rect 119200 19048 120000 19168
rect 119200 17960 120000 18080
rect 0 17416 800 17536
rect 119200 16872 120000 16992
rect 0 15784 800 15904
rect 119200 15784 120000 15904
rect 119200 14696 120000 14816
rect 0 14152 800 14272
rect 119200 13608 120000 13728
rect 0 12520 800 12640
rect 119200 12520 120000 12640
rect 119200 11432 120000 11552
rect 0 10888 800 11008
rect 119200 10344 120000 10464
rect 0 9256 800 9376
rect 119200 9256 120000 9376
rect 119200 8168 120000 8288
rect 0 7624 800 7744
<< obsm3 >>
rect 289 112272 119679 117537
rect 880 111992 119679 112272
rect 289 111728 119679 111992
rect 289 111448 119120 111728
rect 289 110640 119679 111448
rect 880 110360 119120 110640
rect 289 109552 119679 110360
rect 289 109272 119120 109552
rect 289 109008 119679 109272
rect 880 108728 119679 109008
rect 289 108464 119679 108728
rect 289 108184 119120 108464
rect 289 107376 119679 108184
rect 880 107096 119120 107376
rect 289 106288 119679 107096
rect 289 106008 119120 106288
rect 289 105744 119679 106008
rect 880 105464 119679 105744
rect 289 105200 119679 105464
rect 289 104920 119120 105200
rect 289 104112 119679 104920
rect 880 103832 119120 104112
rect 289 103024 119679 103832
rect 289 102744 119120 103024
rect 289 102480 119679 102744
rect 880 102200 119679 102480
rect 289 101936 119679 102200
rect 289 101656 119120 101936
rect 289 100848 119679 101656
rect 880 100568 119120 100848
rect 289 99760 119679 100568
rect 289 99480 119120 99760
rect 289 99216 119679 99480
rect 880 98936 119679 99216
rect 289 98672 119679 98936
rect 289 98392 119120 98672
rect 289 97584 119679 98392
rect 880 97304 119120 97584
rect 289 96496 119679 97304
rect 289 96216 119120 96496
rect 289 95952 119679 96216
rect 880 95672 119679 95952
rect 289 95408 119679 95672
rect 289 95128 119120 95408
rect 289 94320 119679 95128
rect 880 94040 119120 94320
rect 289 93232 119679 94040
rect 289 92952 119120 93232
rect 289 92688 119679 92952
rect 880 92408 119679 92688
rect 289 92144 119679 92408
rect 289 91864 119120 92144
rect 289 91056 119679 91864
rect 880 90776 119120 91056
rect 289 89968 119679 90776
rect 289 89688 119120 89968
rect 289 89424 119679 89688
rect 880 89144 119679 89424
rect 289 88880 119679 89144
rect 289 88600 119120 88880
rect 289 87792 119679 88600
rect 880 87512 119120 87792
rect 289 86704 119679 87512
rect 289 86424 119120 86704
rect 289 86160 119679 86424
rect 880 85880 119679 86160
rect 289 85616 119679 85880
rect 289 85336 119120 85616
rect 289 84528 119679 85336
rect 880 84248 119120 84528
rect 289 83440 119679 84248
rect 289 83160 119120 83440
rect 289 82896 119679 83160
rect 880 82616 119679 82896
rect 289 82352 119679 82616
rect 289 82072 119120 82352
rect 289 81264 119679 82072
rect 880 80984 119120 81264
rect 289 80176 119679 80984
rect 289 79896 119120 80176
rect 289 79632 119679 79896
rect 880 79352 119679 79632
rect 289 79088 119679 79352
rect 289 78808 119120 79088
rect 289 78000 119679 78808
rect 880 77720 119120 78000
rect 289 76912 119679 77720
rect 289 76632 119120 76912
rect 289 76368 119679 76632
rect 880 76088 119679 76368
rect 289 75824 119679 76088
rect 289 75544 119120 75824
rect 289 74736 119679 75544
rect 880 74456 119120 74736
rect 289 73648 119679 74456
rect 289 73368 119120 73648
rect 289 73104 119679 73368
rect 880 72824 119679 73104
rect 289 72560 119679 72824
rect 289 72280 119120 72560
rect 289 71472 119679 72280
rect 880 71192 119120 71472
rect 289 70384 119679 71192
rect 289 70104 119120 70384
rect 289 69840 119679 70104
rect 880 69560 119679 69840
rect 289 69296 119679 69560
rect 289 69016 119120 69296
rect 289 68208 119679 69016
rect 880 67928 119120 68208
rect 289 67120 119679 67928
rect 289 66840 119120 67120
rect 289 66576 119679 66840
rect 880 66296 119679 66576
rect 289 66032 119679 66296
rect 289 65752 119120 66032
rect 289 64944 119679 65752
rect 880 64664 119120 64944
rect 289 63856 119679 64664
rect 289 63576 119120 63856
rect 289 63312 119679 63576
rect 880 63032 119679 63312
rect 289 62768 119679 63032
rect 289 62488 119120 62768
rect 289 61680 119679 62488
rect 880 61400 119120 61680
rect 289 60592 119679 61400
rect 289 60312 119120 60592
rect 289 60048 119679 60312
rect 880 59768 119679 60048
rect 289 59504 119679 59768
rect 289 59224 119120 59504
rect 289 58416 119679 59224
rect 880 58136 119120 58416
rect 289 57328 119679 58136
rect 289 57048 119120 57328
rect 289 56784 119679 57048
rect 880 56504 119679 56784
rect 289 56240 119679 56504
rect 289 55960 119120 56240
rect 289 55152 119679 55960
rect 880 54872 119120 55152
rect 289 54064 119679 54872
rect 289 53784 119120 54064
rect 289 53520 119679 53784
rect 880 53240 119679 53520
rect 289 52976 119679 53240
rect 289 52696 119120 52976
rect 289 51888 119679 52696
rect 880 51608 119120 51888
rect 289 50800 119679 51608
rect 289 50520 119120 50800
rect 289 50256 119679 50520
rect 880 49976 119679 50256
rect 289 49712 119679 49976
rect 289 49432 119120 49712
rect 289 48624 119679 49432
rect 880 48344 119120 48624
rect 289 47536 119679 48344
rect 289 47256 119120 47536
rect 289 46992 119679 47256
rect 880 46712 119679 46992
rect 289 46448 119679 46712
rect 289 46168 119120 46448
rect 289 45360 119679 46168
rect 880 45080 119120 45360
rect 289 44272 119679 45080
rect 289 43992 119120 44272
rect 289 43728 119679 43992
rect 880 43448 119679 43728
rect 289 43184 119679 43448
rect 289 42904 119120 43184
rect 289 42096 119679 42904
rect 880 41816 119120 42096
rect 289 41008 119679 41816
rect 289 40728 119120 41008
rect 289 40464 119679 40728
rect 880 40184 119679 40464
rect 289 39920 119679 40184
rect 289 39640 119120 39920
rect 289 38832 119679 39640
rect 880 38552 119120 38832
rect 289 37744 119679 38552
rect 289 37464 119120 37744
rect 289 37200 119679 37464
rect 880 36920 119679 37200
rect 289 36656 119679 36920
rect 289 36376 119120 36656
rect 289 35568 119679 36376
rect 880 35288 119120 35568
rect 289 34480 119679 35288
rect 289 34200 119120 34480
rect 289 33936 119679 34200
rect 880 33656 119679 33936
rect 289 33392 119679 33656
rect 289 33112 119120 33392
rect 289 32304 119679 33112
rect 880 32024 119120 32304
rect 289 31216 119679 32024
rect 289 30936 119120 31216
rect 289 30672 119679 30936
rect 880 30392 119679 30672
rect 289 30128 119679 30392
rect 289 29848 119120 30128
rect 289 29040 119679 29848
rect 880 28760 119120 29040
rect 289 27952 119679 28760
rect 289 27672 119120 27952
rect 289 27408 119679 27672
rect 880 27128 119679 27408
rect 289 26864 119679 27128
rect 289 26584 119120 26864
rect 289 25776 119679 26584
rect 880 25496 119120 25776
rect 289 24688 119679 25496
rect 289 24408 119120 24688
rect 289 24144 119679 24408
rect 880 23864 119679 24144
rect 289 23600 119679 23864
rect 289 23320 119120 23600
rect 289 22512 119679 23320
rect 880 22232 119120 22512
rect 289 21424 119679 22232
rect 289 21144 119120 21424
rect 289 20880 119679 21144
rect 880 20600 119679 20880
rect 289 20336 119679 20600
rect 289 20056 119120 20336
rect 289 19248 119679 20056
rect 880 18968 119120 19248
rect 289 18160 119679 18968
rect 289 17880 119120 18160
rect 289 17616 119679 17880
rect 880 17336 119679 17616
rect 289 17072 119679 17336
rect 289 16792 119120 17072
rect 289 15984 119679 16792
rect 880 15704 119120 15984
rect 289 14896 119679 15704
rect 289 14616 119120 14896
rect 289 14352 119679 14616
rect 880 14072 119679 14352
rect 289 13808 119679 14072
rect 289 13528 119120 13808
rect 289 12720 119679 13528
rect 880 12440 119120 12720
rect 289 11632 119679 12440
rect 289 11352 119120 11632
rect 289 11088 119679 11352
rect 880 10808 119679 11088
rect 289 10544 119679 10808
rect 289 10264 119120 10544
rect 289 9456 119679 10264
rect 880 9176 119120 9456
rect 289 8368 119679 9176
rect 289 8088 119120 8368
rect 289 7824 119679 8088
rect 880 7544 119679 7824
rect 289 579 119679 7544
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 795 2048 4128 114613
rect 4608 2048 19488 114613
rect 19968 2048 34848 114613
rect 35328 2048 50208 114613
rect 50688 2048 65568 114613
rect 66048 2048 80928 114613
rect 81408 2048 96288 114613
rect 96768 2048 111648 114613
rect 112128 2048 117149 114613
rect 795 579 117149 2048
<< labels >>
rlabel metal2 s 1950 119200 2006 120000 6 clk
port 1 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 dmemreq_addr[0]
port 2 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 dmemreq_addr[10]
port 3 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 dmemreq_addr[11]
port 4 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 dmemreq_addr[12]
port 5 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 dmemreq_addr[13]
port 6 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 dmemreq_addr[14]
port 7 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 dmemreq_addr[15]
port 8 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 dmemreq_addr[16]
port 9 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 dmemreq_addr[17]
port 10 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 dmemreq_addr[18]
port 11 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 dmemreq_addr[19]
port 12 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 dmemreq_addr[1]
port 13 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 dmemreq_addr[20]
port 14 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 dmemreq_addr[21]
port 15 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 dmemreq_addr[22]
port 16 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 dmemreq_addr[23]
port 17 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 dmemreq_addr[24]
port 18 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 dmemreq_addr[25]
port 19 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 dmemreq_addr[26]
port 20 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 dmemreq_addr[27]
port 21 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 dmemreq_addr[28]
port 22 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 dmemreq_addr[29]
port 23 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 dmemreq_addr[2]
port 24 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 dmemreq_addr[30]
port 25 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 dmemreq_addr[31]
port 26 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 dmemreq_addr[3]
port 27 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 dmemreq_addr[4]
port 28 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 dmemreq_addr[5]
port 29 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 dmemreq_addr[6]
port 30 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 dmemreq_addr[7]
port 31 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 dmemreq_addr[8]
port 32 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 dmemreq_addr[9]
port 33 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 dmemreq_type
port 34 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 dmemreq_val
port 35 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 dmemreq_wdata[0]
port 36 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 dmemreq_wdata[10]
port 37 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 dmemreq_wdata[11]
port 38 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 dmemreq_wdata[12]
port 39 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 dmemreq_wdata[13]
port 40 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 dmemreq_wdata[14]
port 41 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 dmemreq_wdata[15]
port 42 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 dmemreq_wdata[16]
port 43 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 dmemreq_wdata[17]
port 44 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 dmemreq_wdata[18]
port 45 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 dmemreq_wdata[19]
port 46 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 dmemreq_wdata[1]
port 47 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 dmemreq_wdata[20]
port 48 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 dmemreq_wdata[21]
port 49 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 dmemreq_wdata[22]
port 50 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 dmemreq_wdata[23]
port 51 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 dmemreq_wdata[24]
port 52 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 dmemreq_wdata[25]
port 53 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 dmemreq_wdata[26]
port 54 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 dmemreq_wdata[27]
port 55 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 dmemreq_wdata[28]
port 56 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 dmemreq_wdata[29]
port 57 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 dmemreq_wdata[2]
port 58 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 dmemreq_wdata[30]
port 59 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 dmemreq_wdata[31]
port 60 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 dmemreq_wdata[3]
port 61 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 dmemreq_wdata[4]
port 62 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 dmemreq_wdata[5]
port 63 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 dmemreq_wdata[6]
port 64 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 dmemreq_wdata[7]
port 65 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 dmemreq_wdata[8]
port 66 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 dmemreq_wdata[9]
port 67 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 dmemresp_rdata[0]
port 68 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 dmemresp_rdata[10]
port 69 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 dmemresp_rdata[11]
port 70 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 dmemresp_rdata[12]
port 71 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 dmemresp_rdata[13]
port 72 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 dmemresp_rdata[14]
port 73 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 dmemresp_rdata[15]
port 74 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 dmemresp_rdata[16]
port 75 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 dmemresp_rdata[17]
port 76 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 dmemresp_rdata[18]
port 77 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 dmemresp_rdata[19]
port 78 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 dmemresp_rdata[1]
port 79 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 dmemresp_rdata[20]
port 80 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 dmemresp_rdata[21]
port 81 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 dmemresp_rdata[22]
port 82 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 dmemresp_rdata[23]
port 83 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 dmemresp_rdata[24]
port 84 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 dmemresp_rdata[25]
port 85 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 dmemresp_rdata[26]
port 86 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 dmemresp_rdata[27]
port 87 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 dmemresp_rdata[28]
port 88 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 dmemresp_rdata[29]
port 89 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 dmemresp_rdata[2]
port 90 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 dmemresp_rdata[30]
port 91 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 dmemresp_rdata[31]
port 92 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 dmemresp_rdata[3]
port 93 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 dmemresp_rdata[4]
port 94 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 dmemresp_rdata[5]
port 95 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 dmemresp_rdata[6]
port 96 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 dmemresp_rdata[7]
port 97 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 dmemresp_rdata[8]
port 98 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 dmemresp_rdata[9]
port 99 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 imemreq_addr[0]
port 100 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 imemreq_addr[10]
port 101 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 imemreq_addr[11]
port 102 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 imemreq_addr[12]
port 103 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 imemreq_addr[13]
port 104 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 imemreq_addr[14]
port 105 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 imemreq_addr[15]
port 106 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 imemreq_addr[16]
port 107 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 imemreq_addr[17]
port 108 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 imemreq_addr[18]
port 109 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 imemreq_addr[19]
port 110 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 imemreq_addr[1]
port 111 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 imemreq_addr[20]
port 112 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 imemreq_addr[21]
port 113 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 imemreq_addr[22]
port 114 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 imemreq_addr[23]
port 115 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 imemreq_addr[24]
port 116 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 imemreq_addr[25]
port 117 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 imemreq_addr[26]
port 118 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 imemreq_addr[27]
port 119 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 imemreq_addr[28]
port 120 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 imemreq_addr[29]
port 121 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 imemreq_addr[2]
port 122 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 imemreq_addr[30]
port 123 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 imemreq_addr[31]
port 124 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 imemreq_addr[3]
port 125 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 imemreq_addr[4]
port 126 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 imemreq_addr[5]
port 127 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 imemreq_addr[6]
port 128 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 imemreq_addr[7]
port 129 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 imemreq_addr[8]
port 130 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 imemreq_addr[9]
port 131 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 imemreq_val
port 132 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 imemresp_data[0]
port 133 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 imemresp_data[10]
port 134 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 imemresp_data[11]
port 135 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 imemresp_data[12]
port 136 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 imemresp_data[13]
port 137 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 imemresp_data[14]
port 138 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 imemresp_data[15]
port 139 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 imemresp_data[16]
port 140 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 imemresp_data[17]
port 141 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 imemresp_data[18]
port 142 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 imemresp_data[19]
port 143 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 imemresp_data[1]
port 144 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 imemresp_data[20]
port 145 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 imemresp_data[21]
port 146 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 imemresp_data[22]
port 147 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 imemresp_data[23]
port 148 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 imemresp_data[24]
port 149 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 imemresp_data[25]
port 150 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 imemresp_data[26]
port 151 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 imemresp_data[27]
port 152 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 imemresp_data[28]
port 153 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 imemresp_data[29]
port 154 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 imemresp_data[2]
port 155 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 imemresp_data[30]
port 156 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 imemresp_data[31]
port 157 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 imemresp_data[3]
port 158 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 imemresp_data[4]
port 159 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 imemresp_data[5]
port 160 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 imemresp_data[6]
port 161 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 imemresp_data[7]
port 162 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 imemresp_data[8]
port 163 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 imemresp_data[9]
port 164 nsew signal input
rlabel metal2 s 4342 119200 4398 120000 6 in0[0]
port 165 nsew signal input
rlabel metal2 s 16302 119200 16358 120000 6 in0[10]
port 166 nsew signal input
rlabel metal2 s 17498 119200 17554 120000 6 in0[11]
port 167 nsew signal input
rlabel metal2 s 18694 119200 18750 120000 6 in0[12]
port 168 nsew signal input
rlabel metal2 s 19890 119200 19946 120000 6 in0[13]
port 169 nsew signal input
rlabel metal2 s 21086 119200 21142 120000 6 in0[14]
port 170 nsew signal input
rlabel metal2 s 22282 119200 22338 120000 6 in0[15]
port 171 nsew signal input
rlabel metal2 s 23478 119200 23534 120000 6 in0[16]
port 172 nsew signal input
rlabel metal2 s 24674 119200 24730 120000 6 in0[17]
port 173 nsew signal input
rlabel metal2 s 25870 119200 25926 120000 6 in0[18]
port 174 nsew signal input
rlabel metal2 s 27066 119200 27122 120000 6 in0[19]
port 175 nsew signal input
rlabel metal2 s 5538 119200 5594 120000 6 in0[1]
port 176 nsew signal input
rlabel metal2 s 28262 119200 28318 120000 6 in0[20]
port 177 nsew signal input
rlabel metal2 s 29458 119200 29514 120000 6 in0[21]
port 178 nsew signal input
rlabel metal2 s 30654 119200 30710 120000 6 in0[22]
port 179 nsew signal input
rlabel metal2 s 31850 119200 31906 120000 6 in0[23]
port 180 nsew signal input
rlabel metal2 s 33046 119200 33102 120000 6 in0[24]
port 181 nsew signal input
rlabel metal2 s 34242 119200 34298 120000 6 in0[25]
port 182 nsew signal input
rlabel metal2 s 35438 119200 35494 120000 6 in0[26]
port 183 nsew signal input
rlabel metal2 s 36634 119200 36690 120000 6 in0[27]
port 184 nsew signal input
rlabel metal2 s 37830 119200 37886 120000 6 in0[28]
port 185 nsew signal input
rlabel metal2 s 39026 119200 39082 120000 6 in0[29]
port 186 nsew signal input
rlabel metal2 s 6734 119200 6790 120000 6 in0[2]
port 187 nsew signal input
rlabel metal2 s 40222 119200 40278 120000 6 in0[30]
port 188 nsew signal input
rlabel metal2 s 41418 119200 41474 120000 6 in0[31]
port 189 nsew signal input
rlabel metal2 s 7930 119200 7986 120000 6 in0[3]
port 190 nsew signal input
rlabel metal2 s 9126 119200 9182 120000 6 in0[4]
port 191 nsew signal input
rlabel metal2 s 10322 119200 10378 120000 6 in0[5]
port 192 nsew signal input
rlabel metal2 s 11518 119200 11574 120000 6 in0[6]
port 193 nsew signal input
rlabel metal2 s 12714 119200 12770 120000 6 in0[7]
port 194 nsew signal input
rlabel metal2 s 13910 119200 13966 120000 6 in0[8]
port 195 nsew signal input
rlabel metal2 s 15106 119200 15162 120000 6 in0[9]
port 196 nsew signal input
rlabel metal2 s 42614 119200 42670 120000 6 in1[0]
port 197 nsew signal input
rlabel metal2 s 54574 119200 54630 120000 6 in1[10]
port 198 nsew signal input
rlabel metal2 s 55770 119200 55826 120000 6 in1[11]
port 199 nsew signal input
rlabel metal2 s 56966 119200 57022 120000 6 in1[12]
port 200 nsew signal input
rlabel metal2 s 58162 119200 58218 120000 6 in1[13]
port 201 nsew signal input
rlabel metal2 s 59358 119200 59414 120000 6 in1[14]
port 202 nsew signal input
rlabel metal2 s 60554 119200 60610 120000 6 in1[15]
port 203 nsew signal input
rlabel metal2 s 61750 119200 61806 120000 6 in1[16]
port 204 nsew signal input
rlabel metal2 s 62946 119200 63002 120000 6 in1[17]
port 205 nsew signal input
rlabel metal2 s 64142 119200 64198 120000 6 in1[18]
port 206 nsew signal input
rlabel metal2 s 65338 119200 65394 120000 6 in1[19]
port 207 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 in1[1]
port 208 nsew signal input
rlabel metal2 s 66534 119200 66590 120000 6 in1[20]
port 209 nsew signal input
rlabel metal2 s 67730 119200 67786 120000 6 in1[21]
port 210 nsew signal input
rlabel metal2 s 68926 119200 68982 120000 6 in1[22]
port 211 nsew signal input
rlabel metal2 s 70122 119200 70178 120000 6 in1[23]
port 212 nsew signal input
rlabel metal2 s 71318 119200 71374 120000 6 in1[24]
port 213 nsew signal input
rlabel metal2 s 72514 119200 72570 120000 6 in1[25]
port 214 nsew signal input
rlabel metal2 s 73710 119200 73766 120000 6 in1[26]
port 215 nsew signal input
rlabel metal2 s 74906 119200 74962 120000 6 in1[27]
port 216 nsew signal input
rlabel metal2 s 76102 119200 76158 120000 6 in1[28]
port 217 nsew signal input
rlabel metal2 s 77298 119200 77354 120000 6 in1[29]
port 218 nsew signal input
rlabel metal2 s 45006 119200 45062 120000 6 in1[2]
port 219 nsew signal input
rlabel metal2 s 78494 119200 78550 120000 6 in1[30]
port 220 nsew signal input
rlabel metal2 s 79690 119200 79746 120000 6 in1[31]
port 221 nsew signal input
rlabel metal2 s 46202 119200 46258 120000 6 in1[3]
port 222 nsew signal input
rlabel metal2 s 47398 119200 47454 120000 6 in1[4]
port 223 nsew signal input
rlabel metal2 s 48594 119200 48650 120000 6 in1[5]
port 224 nsew signal input
rlabel metal2 s 49790 119200 49846 120000 6 in1[6]
port 225 nsew signal input
rlabel metal2 s 50986 119200 51042 120000 6 in1[7]
port 226 nsew signal input
rlabel metal2 s 52182 119200 52238 120000 6 in1[8]
port 227 nsew signal input
rlabel metal2 s 53378 119200 53434 120000 6 in1[9]
port 228 nsew signal input
rlabel metal2 s 80886 119200 80942 120000 6 in2[0]
port 229 nsew signal input
rlabel metal2 s 92846 119200 92902 120000 6 in2[10]
port 230 nsew signal input
rlabel metal2 s 94042 119200 94098 120000 6 in2[11]
port 231 nsew signal input
rlabel metal2 s 95238 119200 95294 120000 6 in2[12]
port 232 nsew signal input
rlabel metal2 s 96434 119200 96490 120000 6 in2[13]
port 233 nsew signal input
rlabel metal2 s 97630 119200 97686 120000 6 in2[14]
port 234 nsew signal input
rlabel metal2 s 98826 119200 98882 120000 6 in2[15]
port 235 nsew signal input
rlabel metal2 s 100022 119200 100078 120000 6 in2[16]
port 236 nsew signal input
rlabel metal2 s 101218 119200 101274 120000 6 in2[17]
port 237 nsew signal input
rlabel metal2 s 102414 119200 102470 120000 6 in2[18]
port 238 nsew signal input
rlabel metal2 s 103610 119200 103666 120000 6 in2[19]
port 239 nsew signal input
rlabel metal2 s 82082 119200 82138 120000 6 in2[1]
port 240 nsew signal input
rlabel metal2 s 104806 119200 104862 120000 6 in2[20]
port 241 nsew signal input
rlabel metal2 s 106002 119200 106058 120000 6 in2[21]
port 242 nsew signal input
rlabel metal2 s 107198 119200 107254 120000 6 in2[22]
port 243 nsew signal input
rlabel metal2 s 108394 119200 108450 120000 6 in2[23]
port 244 nsew signal input
rlabel metal2 s 109590 119200 109646 120000 6 in2[24]
port 245 nsew signal input
rlabel metal2 s 110786 119200 110842 120000 6 in2[25]
port 246 nsew signal input
rlabel metal2 s 111982 119200 112038 120000 6 in2[26]
port 247 nsew signal input
rlabel metal2 s 113178 119200 113234 120000 6 in2[27]
port 248 nsew signal input
rlabel metal2 s 114374 119200 114430 120000 6 in2[28]
port 249 nsew signal input
rlabel metal2 s 115570 119200 115626 120000 6 in2[29]
port 250 nsew signal input
rlabel metal2 s 83278 119200 83334 120000 6 in2[2]
port 251 nsew signal input
rlabel metal2 s 116766 119200 116822 120000 6 in2[30]
port 252 nsew signal input
rlabel metal2 s 117962 119200 118018 120000 6 in2[31]
port 253 nsew signal input
rlabel metal2 s 84474 119200 84530 120000 6 in2[3]
port 254 nsew signal input
rlabel metal2 s 85670 119200 85726 120000 6 in2[4]
port 255 nsew signal input
rlabel metal2 s 86866 119200 86922 120000 6 in2[5]
port 256 nsew signal input
rlabel metal2 s 88062 119200 88118 120000 6 in2[6]
port 257 nsew signal input
rlabel metal2 s 89258 119200 89314 120000 6 in2[7]
port 258 nsew signal input
rlabel metal2 s 90454 119200 90510 120000 6 in2[8]
port 259 nsew signal input
rlabel metal2 s 91650 119200 91706 120000 6 in2[9]
port 260 nsew signal input
rlabel metal3 s 119200 8168 120000 8288 6 out0[0]
port 261 nsew signal output
rlabel metal3 s 119200 19048 120000 19168 6 out0[10]
port 262 nsew signal output
rlabel metal3 s 119200 20136 120000 20256 6 out0[11]
port 263 nsew signal output
rlabel metal3 s 119200 21224 120000 21344 6 out0[12]
port 264 nsew signal output
rlabel metal3 s 119200 22312 120000 22432 6 out0[13]
port 265 nsew signal output
rlabel metal3 s 119200 23400 120000 23520 6 out0[14]
port 266 nsew signal output
rlabel metal3 s 119200 24488 120000 24608 6 out0[15]
port 267 nsew signal output
rlabel metal3 s 119200 25576 120000 25696 6 out0[16]
port 268 nsew signal output
rlabel metal3 s 119200 26664 120000 26784 6 out0[17]
port 269 nsew signal output
rlabel metal3 s 119200 27752 120000 27872 6 out0[18]
port 270 nsew signal output
rlabel metal3 s 119200 28840 120000 28960 6 out0[19]
port 271 nsew signal output
rlabel metal3 s 119200 9256 120000 9376 6 out0[1]
port 272 nsew signal output
rlabel metal3 s 119200 29928 120000 30048 6 out0[20]
port 273 nsew signal output
rlabel metal3 s 119200 31016 120000 31136 6 out0[21]
port 274 nsew signal output
rlabel metal3 s 119200 32104 120000 32224 6 out0[22]
port 275 nsew signal output
rlabel metal3 s 119200 33192 120000 33312 6 out0[23]
port 276 nsew signal output
rlabel metal3 s 119200 34280 120000 34400 6 out0[24]
port 277 nsew signal output
rlabel metal3 s 119200 35368 120000 35488 6 out0[25]
port 278 nsew signal output
rlabel metal3 s 119200 36456 120000 36576 6 out0[26]
port 279 nsew signal output
rlabel metal3 s 119200 37544 120000 37664 6 out0[27]
port 280 nsew signal output
rlabel metal3 s 119200 38632 120000 38752 6 out0[28]
port 281 nsew signal output
rlabel metal3 s 119200 39720 120000 39840 6 out0[29]
port 282 nsew signal output
rlabel metal3 s 119200 10344 120000 10464 6 out0[2]
port 283 nsew signal output
rlabel metal3 s 119200 40808 120000 40928 6 out0[30]
port 284 nsew signal output
rlabel metal3 s 119200 41896 120000 42016 6 out0[31]
port 285 nsew signal output
rlabel metal3 s 119200 11432 120000 11552 6 out0[3]
port 286 nsew signal output
rlabel metal3 s 119200 12520 120000 12640 6 out0[4]
port 287 nsew signal output
rlabel metal3 s 119200 13608 120000 13728 6 out0[5]
port 288 nsew signal output
rlabel metal3 s 119200 14696 120000 14816 6 out0[6]
port 289 nsew signal output
rlabel metal3 s 119200 15784 120000 15904 6 out0[7]
port 290 nsew signal output
rlabel metal3 s 119200 16872 120000 16992 6 out0[8]
port 291 nsew signal output
rlabel metal3 s 119200 17960 120000 18080 6 out0[9]
port 292 nsew signal output
rlabel metal3 s 119200 42984 120000 43104 6 out1[0]
port 293 nsew signal output
rlabel metal3 s 119200 53864 120000 53984 6 out1[10]
port 294 nsew signal output
rlabel metal3 s 119200 54952 120000 55072 6 out1[11]
port 295 nsew signal output
rlabel metal3 s 119200 56040 120000 56160 6 out1[12]
port 296 nsew signal output
rlabel metal3 s 119200 57128 120000 57248 6 out1[13]
port 297 nsew signal output
rlabel metal3 s 119200 58216 120000 58336 6 out1[14]
port 298 nsew signal output
rlabel metal3 s 119200 59304 120000 59424 6 out1[15]
port 299 nsew signal output
rlabel metal3 s 119200 60392 120000 60512 6 out1[16]
port 300 nsew signal output
rlabel metal3 s 119200 61480 120000 61600 6 out1[17]
port 301 nsew signal output
rlabel metal3 s 119200 62568 120000 62688 6 out1[18]
port 302 nsew signal output
rlabel metal3 s 119200 63656 120000 63776 6 out1[19]
port 303 nsew signal output
rlabel metal3 s 119200 44072 120000 44192 6 out1[1]
port 304 nsew signal output
rlabel metal3 s 119200 64744 120000 64864 6 out1[20]
port 305 nsew signal output
rlabel metal3 s 119200 65832 120000 65952 6 out1[21]
port 306 nsew signal output
rlabel metal3 s 119200 66920 120000 67040 6 out1[22]
port 307 nsew signal output
rlabel metal3 s 119200 68008 120000 68128 6 out1[23]
port 308 nsew signal output
rlabel metal3 s 119200 69096 120000 69216 6 out1[24]
port 309 nsew signal output
rlabel metal3 s 119200 70184 120000 70304 6 out1[25]
port 310 nsew signal output
rlabel metal3 s 119200 71272 120000 71392 6 out1[26]
port 311 nsew signal output
rlabel metal3 s 119200 72360 120000 72480 6 out1[27]
port 312 nsew signal output
rlabel metal3 s 119200 73448 120000 73568 6 out1[28]
port 313 nsew signal output
rlabel metal3 s 119200 74536 120000 74656 6 out1[29]
port 314 nsew signal output
rlabel metal3 s 119200 45160 120000 45280 6 out1[2]
port 315 nsew signal output
rlabel metal3 s 119200 75624 120000 75744 6 out1[30]
port 316 nsew signal output
rlabel metal3 s 119200 76712 120000 76832 6 out1[31]
port 317 nsew signal output
rlabel metal3 s 119200 46248 120000 46368 6 out1[3]
port 318 nsew signal output
rlabel metal3 s 119200 47336 120000 47456 6 out1[4]
port 319 nsew signal output
rlabel metal3 s 119200 48424 120000 48544 6 out1[5]
port 320 nsew signal output
rlabel metal3 s 119200 49512 120000 49632 6 out1[6]
port 321 nsew signal output
rlabel metal3 s 119200 50600 120000 50720 6 out1[7]
port 322 nsew signal output
rlabel metal3 s 119200 51688 120000 51808 6 out1[8]
port 323 nsew signal output
rlabel metal3 s 119200 52776 120000 52896 6 out1[9]
port 324 nsew signal output
rlabel metal3 s 119200 77800 120000 77920 6 out2[0]
port 325 nsew signal output
rlabel metal3 s 119200 88680 120000 88800 6 out2[10]
port 326 nsew signal output
rlabel metal3 s 119200 89768 120000 89888 6 out2[11]
port 327 nsew signal output
rlabel metal3 s 119200 90856 120000 90976 6 out2[12]
port 328 nsew signal output
rlabel metal3 s 119200 91944 120000 92064 6 out2[13]
port 329 nsew signal output
rlabel metal3 s 119200 93032 120000 93152 6 out2[14]
port 330 nsew signal output
rlabel metal3 s 119200 94120 120000 94240 6 out2[15]
port 331 nsew signal output
rlabel metal3 s 119200 95208 120000 95328 6 out2[16]
port 332 nsew signal output
rlabel metal3 s 119200 96296 120000 96416 6 out2[17]
port 333 nsew signal output
rlabel metal3 s 119200 97384 120000 97504 6 out2[18]
port 334 nsew signal output
rlabel metal3 s 119200 98472 120000 98592 6 out2[19]
port 335 nsew signal output
rlabel metal3 s 119200 78888 120000 79008 6 out2[1]
port 336 nsew signal output
rlabel metal3 s 119200 99560 120000 99680 6 out2[20]
port 337 nsew signal output
rlabel metal3 s 119200 100648 120000 100768 6 out2[21]
port 338 nsew signal output
rlabel metal3 s 119200 101736 120000 101856 6 out2[22]
port 339 nsew signal output
rlabel metal3 s 119200 102824 120000 102944 6 out2[23]
port 340 nsew signal output
rlabel metal3 s 119200 103912 120000 104032 6 out2[24]
port 341 nsew signal output
rlabel metal3 s 119200 105000 120000 105120 6 out2[25]
port 342 nsew signal output
rlabel metal3 s 119200 106088 120000 106208 6 out2[26]
port 343 nsew signal output
rlabel metal3 s 119200 107176 120000 107296 6 out2[27]
port 344 nsew signal output
rlabel metal3 s 119200 108264 120000 108384 6 out2[28]
port 345 nsew signal output
rlabel metal3 s 119200 109352 120000 109472 6 out2[29]
port 346 nsew signal output
rlabel metal3 s 119200 79976 120000 80096 6 out2[2]
port 347 nsew signal output
rlabel metal3 s 119200 110440 120000 110560 6 out2[30]
port 348 nsew signal output
rlabel metal3 s 119200 111528 120000 111648 6 out2[31]
port 349 nsew signal output
rlabel metal3 s 119200 81064 120000 81184 6 out2[3]
port 350 nsew signal output
rlabel metal3 s 119200 82152 120000 82272 6 out2[4]
port 351 nsew signal output
rlabel metal3 s 119200 83240 120000 83360 6 out2[5]
port 352 nsew signal output
rlabel metal3 s 119200 84328 120000 84448 6 out2[6]
port 353 nsew signal output
rlabel metal3 s 119200 85416 120000 85536 6 out2[7]
port 354 nsew signal output
rlabel metal3 s 119200 86504 120000 86624 6 out2[8]
port 355 nsew signal output
rlabel metal3 s 119200 87592 120000 87712 6 out2[9]
port 356 nsew signal output
rlabel metal2 s 3146 119200 3202 120000 6 rst
port 357 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 358 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 358 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 358 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 358 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 359 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 359 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 359 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 359 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 41493950
string GDS_FILE /home/js2992/c2s2/tinyrv1/caravel/openlane/Proc/runs/25_02_25_22_09/results/signoff/Proc.magic.gds
string GDS_START 1270678
<< end >>


`ifndef PROCCTRL_V
`define PROCCTRL_V

module ProcCtrl
(

);


endmodule

`endif
* NGSPICE file created from Proc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt Proc clk dmemreq_addr[0] dmemreq_addr[10] dmemreq_addr[11] dmemreq_addr[12]
+ dmemreq_addr[13] dmemreq_addr[14] dmemreq_addr[15] dmemreq_addr[16] dmemreq_addr[17]
+ dmemreq_addr[18] dmemreq_addr[19] dmemreq_addr[1] dmemreq_addr[20] dmemreq_addr[21]
+ dmemreq_addr[22] dmemreq_addr[23] dmemreq_addr[24] dmemreq_addr[25] dmemreq_addr[26]
+ dmemreq_addr[27] dmemreq_addr[28] dmemreq_addr[29] dmemreq_addr[2] dmemreq_addr[30]
+ dmemreq_addr[31] dmemreq_addr[3] dmemreq_addr[4] dmemreq_addr[5] dmemreq_addr[6]
+ dmemreq_addr[7] dmemreq_addr[8] dmemreq_addr[9] dmemreq_type dmemreq_val dmemreq_wdata[0]
+ dmemreq_wdata[10] dmemreq_wdata[11] dmemreq_wdata[12] dmemreq_wdata[13] dmemreq_wdata[14]
+ dmemreq_wdata[15] dmemreq_wdata[16] dmemreq_wdata[17] dmemreq_wdata[18] dmemreq_wdata[19]
+ dmemreq_wdata[1] dmemreq_wdata[20] dmemreq_wdata[21] dmemreq_wdata[22] dmemreq_wdata[23]
+ dmemreq_wdata[24] dmemreq_wdata[25] dmemreq_wdata[26] dmemreq_wdata[27] dmemreq_wdata[28]
+ dmemreq_wdata[29] dmemreq_wdata[2] dmemreq_wdata[30] dmemreq_wdata[31] dmemreq_wdata[3]
+ dmemreq_wdata[4] dmemreq_wdata[5] dmemreq_wdata[6] dmemreq_wdata[7] dmemreq_wdata[8]
+ dmemreq_wdata[9] dmemresp_rdata[0] dmemresp_rdata[10] dmemresp_rdata[11] dmemresp_rdata[12]
+ dmemresp_rdata[13] dmemresp_rdata[14] dmemresp_rdata[15] dmemresp_rdata[16] dmemresp_rdata[17]
+ dmemresp_rdata[18] dmemresp_rdata[19] dmemresp_rdata[1] dmemresp_rdata[20] dmemresp_rdata[21]
+ dmemresp_rdata[22] dmemresp_rdata[23] dmemresp_rdata[24] dmemresp_rdata[25] dmemresp_rdata[26]
+ dmemresp_rdata[27] dmemresp_rdata[28] dmemresp_rdata[29] dmemresp_rdata[2] dmemresp_rdata[30]
+ dmemresp_rdata[31] dmemresp_rdata[3] dmemresp_rdata[4] dmemresp_rdata[5] dmemresp_rdata[6]
+ dmemresp_rdata[7] dmemresp_rdata[8] dmemresp_rdata[9] imemreq_addr[0] imemreq_addr[10]
+ imemreq_addr[11] imemreq_addr[12] imemreq_addr[13] imemreq_addr[14] imemreq_addr[15]
+ imemreq_addr[16] imemreq_addr[17] imemreq_addr[18] imemreq_addr[19] imemreq_addr[1]
+ imemreq_addr[20] imemreq_addr[21] imemreq_addr[22] imemreq_addr[23] imemreq_addr[24]
+ imemreq_addr[25] imemreq_addr[26] imemreq_addr[27] imemreq_addr[28] imemreq_addr[29]
+ imemreq_addr[2] imemreq_addr[30] imemreq_addr[31] imemreq_addr[3] imemreq_addr[4]
+ imemreq_addr[5] imemreq_addr[6] imemreq_addr[7] imemreq_addr[8] imemreq_addr[9]
+ imemreq_val imemresp_data[0] imemresp_data[10] imemresp_data[11] imemresp_data[12]
+ imemresp_data[13] imemresp_data[14] imemresp_data[15] imemresp_data[16] imemresp_data[17]
+ imemresp_data[18] imemresp_data[19] imemresp_data[1] imemresp_data[20] imemresp_data[21]
+ imemresp_data[22] imemresp_data[23] imemresp_data[24] imemresp_data[25] imemresp_data[26]
+ imemresp_data[27] imemresp_data[28] imemresp_data[29] imemresp_data[2] imemresp_data[30]
+ imemresp_data[31] imemresp_data[3] imemresp_data[4] imemresp_data[5] imemresp_data[6]
+ imemresp_data[7] imemresp_data[8] imemresp_data[9] in0[0] in0[10] in0[11] in0[12]
+ in0[13] in0[14] in0[15] in0[16] in0[17] in0[18] in0[19] in0[1] in0[20] in0[21] in0[22]
+ in0[23] in0[24] in0[25] in0[26] in0[27] in0[28] in0[29] in0[2] in0[30] in0[31] in0[3]
+ in0[4] in0[5] in0[6] in0[7] in0[8] in0[9] in1[0] in1[10] in1[11] in1[12] in1[13]
+ in1[14] in1[15] in1[16] in1[17] in1[18] in1[19] in1[1] in1[20] in1[21] in1[22] in1[23]
+ in1[24] in1[25] in1[26] in1[27] in1[28] in1[29] in1[2] in1[30] in1[31] in1[3] in1[4]
+ in1[5] in1[6] in1[7] in1[8] in1[9] in2[0] in2[10] in2[11] in2[12] in2[13] in2[14]
+ in2[15] in2[16] in2[17] in2[18] in2[19] in2[1] in2[20] in2[21] in2[22] in2[23] in2[24]
+ in2[25] in2[26] in2[27] in2[28] in2[29] in2[2] in2[30] in2[31] in2[3] in2[4] in2[5]
+ in2[6] in2[7] in2[8] in2[9] out0[0] out0[10] out0[11] out0[12] out0[13] out0[14]
+ out0[15] out0[16] out0[17] out0[18] out0[19] out0[1] out0[20] out0[21] out0[22]
+ out0[23] out0[24] out0[25] out0[26] out0[27] out0[28] out0[29] out0[2] out0[30]
+ out0[31] out0[3] out0[4] out0[5] out0[6] out0[7] out0[8] out0[9] out1[0] out1[10]
+ out1[11] out1[12] out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19]
+ out1[1] out1[20] out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27]
+ out1[28] out1[29] out1[2] out1[30] out1[31] out1[3] out1[4] out1[5] out1[6] out1[7]
+ out1[8] out1[9] out2[0] out2[10] out2[11] out2[12] out2[13] out2[14] out2[15] out2[16]
+ out2[17] out2[18] out2[19] out2[1] out2[20] out2[21] out2[22] out2[23] out2[24]
+ out2[25] out2[26] out2[27] out2[28] out2[29] out2[2] out2[30] out2[31] out2[3] out2[4]
+ out2[5] out2[6] out2[7] out2[8] out2[9] rst vccd1 vssd1
XANTENNA__12202__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07534__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ _08621_/B _08621_/C _08621_/A vssd1 vssd1 vccd1 vccd1 _08622_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08553_ _08981_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08553_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07504_ hold1007/X _13743_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07504_/X sky130_fd_sc_hd__mux2_1
X_08484_ _08483_/A _08483_/B _08483_/C vssd1 vssd1 vccd1 vccd1 _08485_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_159_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07435_ _08849_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14065_/D sky130_fd_sc_hd__and2_1
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12665__S _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout427_A _11829_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07759__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ _15349_/Q _14062_/Q vssd1 vssd1 vccd1 vccd1 _07366_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10693__B _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12594__A1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _09941_/A _09105_/B vssd1 vssd1 vccd1 vccd1 _09105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07297_ _11620_/B _14964_/Q vssd1 vssd1 vccd1 vccd1 _07297_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08262__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ _09164_/A _09979_/C vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout796_A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold340 hold340/A vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10357__B1 _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 hold351/A vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07494__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold362 hold362/A vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 hold373/A vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 hold384/A vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold395 hold395/A vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _12460_/S vssd1 vssd1 vccd1 vccd1 _12459_/S sky130_fd_sc_hd__buf_6
XANTENNA__08970__B1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 _12791_/S vssd1 vssd1 vccd1 vccd1 _12735_/S sky130_fd_sc_hd__buf_8
XANTENNA__10109__B1 _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _11507_/A _09935_/X _09937_/X vssd1 vssd1 vccd1 vccd1 _09938_/Y sky130_fd_sc_hd__o21ai_1
Xfanout842 _14488_/Q vssd1 vssd1 vccd1 vccd1 _12964_/S0 sky130_fd_sc_hd__buf_6
Xfanout853 _13622_/C1 vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__buf_4
XFILLER_0_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout864 _13404_/A vssd1 vssd1 vccd1 vccd1 _13397_/A sky130_fd_sc_hd__clkbuf_4
Xfanout875 _13501_/A vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__buf_4
XFILLER_0_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout886 _13168_/A vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__clkbuf_4
X_09869_ _09869_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__and3_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 _13205_/X vssd1 vssd1 vccd1 vccd1 _15069_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11744__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 _14725_/Q vssd1 vssd1 vccd1 vccd1 hold1051/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1062 _07628_/X vssd1 vssd1 vccd1 vccd1 _14251_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ _13655_/A1 hold1399/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11900_/X sky130_fd_sc_hd__mux2_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1073 _13972_/Q vssd1 vssd1 vccd1 vccd1 hold1073/X sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _13080_/A1 _12879_/X _12877_/X vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__a21oi_4
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 _07494_/X vssd1 vssd1 vccd1 vccd1 _14122_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _14358_/Q vssd1 vssd1 vccd1 vccd1 hold1095/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_202 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ hold853/X hold2816/X _11845_/S vssd1 vssd1 vccd1 vccd1 hold854/A sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09278__A1 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_224 _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__B _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07242__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ _15415_/CLK hold984/X vssd1 vssd1 vccd1 vccd1 hold983/A sky130_fd_sc_hd__dfxtp_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09373__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _13715_/A1 hold1641/X _11762_/S vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__mux2_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13501_ _13501_/A hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__and2_1
XFILLER_0_138_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10713_ _10713_/A _10713_/B _10713_/C vssd1 vssd1 vccd1 vccd1 _10713_/Y sky130_fd_sc_hd__nor3_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _15415_/CLK _14481_/D vssd1 vssd1 vccd1 vccd1 _14481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ input49/X _13648_/B vssd1 vssd1 vccd1 vccd1 _11693_/X sky130_fd_sc_hd__or2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13260__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12034__A0 hold2439/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07669__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ _08851_/A _12273_/B _13440_/S vssd1 vssd1 vccd1 vccd1 _13433_/B sky130_fd_sc_hd__mux2_1
X_10644_ _11606_/A _11536_/A _10827_/C _11542_/A vssd1 vssd1 vccd1 vccd1 _10646_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11388__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13369_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _15154_/D sky130_fd_sc_hd__nor2_1
X_10575_ _13749_/A _13456_/B _10574_/X vssd1 vssd1 vccd1 vccd1 _10575_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08073__B _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ _15116_/CLK _15102_/D vssd1 vssd1 vccd1 vccd1 _15102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _15390_/Q hold439/A _14685_/Q _14749_/Q _12365_/S0 _12343_/A vssd1 vssd1
+ vccd1 vccd1 _12314_/X sky130_fd_sc_hd__mux4_1
X_13294_ input137/X fanout5/X fanout3/X input105/X vssd1 vssd1 vccd1 vccd1 _13294_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10108__B _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13534__A0 _15068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output179_A _15190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11919__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ _15196_/CLK _15033_/D vssd1 vssd1 vccd1 vccd1 _15033_/Q sky130_fd_sc_hd__dfxtp_1
X_12245_ _12247_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _12245_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12176_ _14899_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12176_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12323__B _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11560__A2 _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07417__B _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _11509_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11127_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_208_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12196__S0 _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11058_ _11620_/A _11542_/B _10821_/X _10822_/X _11378_/D vssd1 vssd1 vccd1 vccd1
+ _11063_/A sky130_fd_sc_hd__a32o_1
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07516__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11654__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10009_ _10115_/B _10010_/B _10010_/C _10010_/D vssd1 vssd1 vccd1 vccd1 _10011_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14817_ _14840_/CLK _14817_/D vssd1 vssd1 vccd1 vccd1 _14817_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13154__B _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12499__S1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ _15387_/CLK hold992/X vssd1 vssd1 vccd1 vccd1 hold991/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10823__A1 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12485__S _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14679_ _15453_/CLK _14679_/D vssd1 vssd1 vccd1 vccd1 _14679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07220_ hold262/A _07855_/A _07218_/X _07856_/B vssd1 vssd1 vccd1 vccd1 _07221_/A
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ _13652_/A1 hold1943/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07151_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_171_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2559_A _12276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12671__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07082_ _13718_/A1 hold1591/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07082_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12328__A1 _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold2726_A _15178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10339__B1 _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12879__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12423__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11000__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11000__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09526__C _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__A3 _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07984_ _13866_/Q _13994_/Q hold809/A hold929/A _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07984_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_199_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09723_ _10115_/B _09724_/C _09724_/D _10115_/A vssd1 vssd1 vccd1 vccd1 _09726_/C
+ sky130_fd_sc_hd__a22o_1
X_06935_ _06935_/A vssd1 vssd1 vccd1 vccd1 _06935_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10969__A _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07507__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout377_A _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _13704_/A1 _11514_/A2 _11514_/B1 _13192_/B _09652_/Y vssd1 vssd1 vccd1 vccd1
+ _09654_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_78_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08605_ _08926_/A _08702_/B _08604_/C _08699_/A vssd1 vssd1 vccd1 vccd1 _08606_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _09585_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _09587_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_49_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout544_A _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08536_ _08536_/A _08536_/B vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13461__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08467_ _13661_/A1 _12260_/A2 _12259_/A1 _13182_/B _08465_/Y vssd1 vssd1 vccd1 vccd1
+ _08467_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout809_A _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__A0 hold2602/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07418_ hold19/X _07473_/B vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__and2_1
X_08398_ _08397_/B _08397_/C _08397_/A vssd1 vssd1 vccd1 vccd1 _08400_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_46_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ _07353_/D _15330_/Q vssd1 vssd1 vccd1 vccd1 _07360_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_163_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _10360_/A _10524_/B _10360_/C vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11739__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09019_ _09146_/A _09019_/B vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__and2_1
XFILLER_0_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10291_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12414__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ hold2509/X hold2674/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10425__S0 _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13239__B _15352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_151_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout650 _08677_/A vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_31_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout661 hold2742/X vssd1 vssd1 vccd1 vccd1 _13679_/A1 sky130_fd_sc_hd__buf_4
Xfanout672 _15060_/Q vssd1 vssd1 vccd1 vccd1 _13740_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_205_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout683 _15055_/Q vssd1 vssd1 vccd1 vccd1 _13735_/A1 sky130_fd_sc_hd__buf_4
X_13981_ _14612_/CLK _13981_/D vssd1 vssd1 vccd1 vccd1 _13981_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10879__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout694 _13729_/A1 vssd1 vssd1 vccd1 vccd1 _13663_/A1 sky130_fd_sc_hd__buf_4
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12932_ _13171_/A _12932_/B vssd1 vssd1 vccd1 vccd1 _14965_/D sky130_fd_sc_hd__nor2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_166_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07253__A _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12917_/B1 _12858_/X _12862_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12870_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11058__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/CLK hold698/X vssd1 vssd1 vccd1 vccd1 hold697/A sky130_fd_sc_hd__dfxtp_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ hold351/X _13668_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold352/A sky130_fd_sc_hd__mux2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11058__B2 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12255__B1 _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12794_ _12844_/A1 _12789_/X _12793_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12795_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14533_ _15435_/CLK _14533_/D vssd1 vssd1 vccd1 vccd1 _14533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _13698_/A1 hold653/X _11745_/S vssd1 vssd1 vccd1 vccd1 hold654/A sky130_fd_sc_hd__mux2_1
XFILLER_0_200_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14464_ _15398_/CLK _14464_/D vssd1 vssd1 vccd1 vccd1 _14464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11676_ _13740_/A1 hold2171/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_165_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ _08038_/A _13466_/A _13414_/Y _13178_/A vssd1 vssd1 vccd1 vccd1 _15201_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10627_ _10627_/A _10795_/A _10627_/C vssd1 vssd1 vccd1 vccd1 _10795_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14395_ _15360_/CLK _14395_/D vssd1 vssd1 vccd1 vccd1 _14395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ _13360_/A _13346_/B vssd1 vssd1 vccd1 vccd1 _15137_/D sky130_fd_sc_hd__nor2_1
X_10558_ _10558_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10560_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07985__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ input67/X fanout1/X _13276_/X vssd1 vssd1 vccd1 vccd1 _13278_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12334__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ _10489_/A _10652_/B _10489_/C vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_122_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10780__C _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15016_ _15179_/CLK _15016_/D vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__dfxtp_1
X_12228_ hold251/A hold743/A hold907/A _13959_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12229_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13149__B _13149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12730__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ hold2538/X _12195_/A2 _12158_/X _13491_/A vssd1 vssd1 vccd1 vccd1 _12159_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1809 _14647_/Q vssd1 vssd1 vccd1 vccd1 hold1809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09643__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13165__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _10426_/A _09370_/B vssd1 vssd1 vccd1 vccd1 _09370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09111__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08321_ _08320_/A _08320_/B _08413_/A _08320_/D vssd1 vssd1 vccd1 vccd1 _08322_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08252_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_157_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08870__C1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ hold617/X _13671_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold618/A sky130_fd_sc_hd__mux2_1
XANTENNA__07102__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _09918_/A _08176_/Y _13348_/B _08256_/A _08182_/Y vssd1 vssd1 vccd1 vccd1
+ _08183_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11226__A2_N _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07134_ _13735_/A1 hold2229/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07134_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07065_ _13703_/A1 hold1287/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07065_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput220 _14201_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[31] sky130_fd_sc_hd__buf_12
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08441__B _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput231 _14436_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[12] sky130_fd_sc_hd__buf_12
XFILLER_0_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput242 _14446_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[22] sky130_fd_sc_hd__buf_12
XFILLER_0_140_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput253 _14427_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[3] sky130_fd_sc_hd__buf_12
Xoutput264 _14890_/Q vssd1 vssd1 vccd1 vccd1 out0[13] sky130_fd_sc_hd__buf_12
XFILLER_0_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput275 _14900_/Q vssd1 vssd1 vccd1 vccd1 out0[23] sky130_fd_sc_hd__buf_12
XANTENNA_fanout494_A _06944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput286 _14881_/Q vssd1 vssd1 vccd1 vccd1 out0[4] sky130_fd_sc_hd__buf_12
Xoutput297 _14859_/Q vssd1 vssd1 vccd1 vccd1 out1[14] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07772__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ hold2788/X _07966_/Y _12256_/A vssd1 vssd1 vccd1 vccd1 _07967_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_199_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09706_ _09706_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11288__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06918_ _06918_/A vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__inv_2
X_07898_ _12221_/B _07887_/Y _07897_/X vssd1 vssd1 vccd1 vccd1 _13376_/B sky130_fd_sc_hd__a21o_4
X_09637_ hold377/A _15281_/Q hold307/A _14382_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09637_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13029__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09568_ _09568_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12788__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08519_ _08519_/A _08519_/B vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _09497_/Y _09780_/B _07390_/A vssd1 vssd1 vccd1 vccd1 _09499_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12883__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ _11366_/X _11368_/Y _11340_/A _15227_/Q vssd1 vssd1 vccd1 vccd1 _11532_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout4_A fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11042__B _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09405__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11461_ _11461_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08208__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _13479_/A _13200_/B vssd1 vssd1 vccd1 vccd1 _15065_/D sky130_fd_sc_hd__and2_1
X_10412_ _11104_/A _12284_/B _10408_/Y _10411_/X vssd1 vssd1 vccd1 vccd1 _10412_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ _11392_/A _11392_/B _11392_/C vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__nand3_2
X_14180_ _15179_/CLK _14180_/D vssd1 vssd1 vccd1 vccd1 _14180_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09500__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ _13495_/A hold117/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__and2_1
X_10343_ _10343_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10345_/B sky130_fd_sc_hd__or2_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09169__B1 _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07248__A _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12399__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _10293_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10294_/A sky130_fd_sc_hd__nand2_1
X_13062_ _13068_/A1 _13059_/X _13061_/X vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12712__A1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13684__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _12063_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _14819_/D sky130_fd_sc_hd__and2_1
XFILLER_0_79_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07682__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout480 _06959_/X vssd1 vssd1 vccd1 vccd1 _12253_/S sky130_fd_sc_hd__buf_6
XFILLER_0_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout491 _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12675_/S1 sky130_fd_sc_hd__buf_8
X_13964_ _14595_/CLK _13964_/D vssd1 vssd1 vccd1 vccd1 _13964_/Q sky130_fd_sc_hd__dfxtp_1
X_12915_ hold897/A _14130_/Q _12915_/S vssd1 vssd1 vccd1 vccd1 _12915_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12571__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13895_ _15428_/CLK _13895_/D vssd1 vssd1 vccd1 vccd1 _13895_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11932__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12846_ hold447/A _15282_/Q _15090_/Q _14383_/Q _12915_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12846_/X sky130_fd_sc_hd__mux4_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__A1 _13392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _13102_/A _12777_/B _12777_/C vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__B _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11233__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12874__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14516_ _15408_/CLK hold650/X vssd1 vssd1 vccd1 vccd1 hold649/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ hold385/X _15068_/Q _11728_/S vssd1 vssd1 vccd1 vccd1 hold386/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14447_ _15423_/CLK _14447_/D vssd1 vssd1 vccd1 vccd1 _14447_/Q sky130_fd_sc_hd__dfxtp_1
X_11659_ _13690_/A1 hold2241/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10006__A2 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__A1 _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14378_ _14472_/CLK _14378_/D vssd1 vssd1 vccd1 vccd1 _14378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold906 hold906/A vssd1 vssd1 vccd1 vccd1 hold906/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold917 hold917/A vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _13338_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _15129_/D sky130_fd_sc_hd__nor2_1
Xhold928 hold928/A vssd1 vssd1 vccd1 vccd1 hold928/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold939 hold939/A vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__B1 _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2307 hold2835/X vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ _08065_/A _08867_/X _08869_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08871_/B
+ sky130_fd_sc_hd__o211a_1
Xhold2318 _07452_/X vssd1 vssd1 vccd1 vccd1 _14082_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2329 _11488_/X vssd1 vssd1 vccd1 vccd1 hold2329/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07592__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09580__B1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1606 _11973_/X vssd1 vssd1 vccd1 vccd1 _14792_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07821_ _14783_/Q _14495_/Q _07822_/S vssd1 vssd1 vccd1 vccd1 _07821_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1617 _14657_/Q vssd1 vssd1 vccd1 vccd1 hold1617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 _07167_/X vssd1 vssd1 vccd1 vccd1 _13975_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1639 _13982_/Q vssd1 vssd1 vccd1 vccd1 hold1639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12467__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _13690_/A1 hold1713/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07752_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08135__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07683_ hold1587/X _13656_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 _07683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11842__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _09420_/B _09420_/C _09420_/A vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12314__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _15150_/Q _09925_/A2 _13570_/B vssd1 vssd1 vccd1 vccd1 _09353_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09635__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08438__A2 _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ _08776_/B _09026_/B _09138_/A _10507_/A vssd1 vssd1 vccd1 vccd1 _08306_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11143__A _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09284_ _10166_/A _10338_/B _09860_/B _09676_/D vssd1 vssd1 vccd1 vccd1 _09285_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_145_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08235_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08326_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10982__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout507_A _06926_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07767__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08166_ _08097_/B _08098_/Y _08097_/A vssd1 vssd1 vccd1 vccd1 _08166_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_0_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08452__A _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07117_ _13718_/A1 hold1717/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07117_/X sky130_fd_sc_hd__mux2_1
X_08097_ _08097_/A _08097_/B vssd1 vssd1 vccd1 vccd1 _08097_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07048_ _13653_/A1 hold2049/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07048_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12155__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12702__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09797__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2830 _15319_/Q vssd1 vssd1 vccd1 vccd1 hold2830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2841 _15297_/Q vssd1 vssd1 vccd1 vccd1 hold2841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2852 _15350_/Q vssd1 vssd1 vccd1 vccd1 hold2852/X sky130_fd_sc_hd__dlygate4sd3_1
X_08999_ _11580_/A _09846_/B _09724_/C vssd1 vssd1 vccd1 vccd1 _09124_/B sky130_fd_sc_hd__and3_1
XFILLER_0_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13009__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07007__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ _11578_/A _14968_/Q _14969_/Q _11580_/A vssd1 vssd1 vccd1 vccd1 _10961_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09874__A1 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11752__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ _12696_/X _12697_/X _12699_/X _12698_/X _12700_/S0 _12700_/S1 vssd1 vssd1
+ vccd1 vccd1 _12701_/B sky130_fd_sc_hd__mux4_1
X_13680_ hold1331/X _13680_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__mux2_1
X_10892_ _10889_/Y _10890_/X _10707_/Y _10709_/X vssd1 vssd1 vccd1 vccd1 _10893_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12631_ _13106_/A1 _13152_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12632_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_39_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _15425_/CLK _15350_/D vssd1 vssd1 vccd1 vccd1 _15350_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10236__A2 _13452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ _12368_/A _12559_/X _12561_/X vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ _15072_/CLK hold404/X vssd1 vssd1 vccd1 vccd1 hold403/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11513_ hold2769/X input25/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13203_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13679__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ _15378_/CLK _15281_/D vssd1 vssd1 vccd1 vccd1 _15281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12493_ _12599_/S1 _12490_/X _12492_/X vssd1 vssd1 vccd1 vccd1 _12493_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12608__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14232_ _14958_/CLK hold824/X vssd1 vssd1 vccd1 vccd1 hold823/A sky130_fd_sc_hd__dfxtp_1
X_11444_ _11443_/B _11443_/C _11443_/A vssd1 vssd1 vccd1 vccd1 _11445_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12394__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14163_ _15415_/CLK hold478/X vssd1 vssd1 vccd1 vccd1 hold477/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08601__A2 _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11375_ _11620_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10095__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ _13491_/A hold51/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__and2_1
XFILLER_0_81_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10326_ _10326_/A _10326_/B _10326_/C vssd1 vssd1 vccd1 vccd1 _10328_/B sky130_fd_sc_hd__and3_2
X_14094_ _14973_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 _14094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09237__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13033__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ _13045_/A _13045_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _13052_/B sky130_fd_sc_hd__or3b_1
Xclkbuf_4_2__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_2__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _11320_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09562__B1 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10188_ _10185_/X _10186_/Y _10019_/D _10020_/B vssd1 vssd1 vccd1 vccd1 _10189_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10132__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14996_ _15004_/CLK hold118/X vssd1 vssd1 vccd1 vccd1 _14996_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08117__A1 _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13947_ _15448_/CLK _13947_/D vssd1 vssd1 vccd1 vccd1 _13947_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11121__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11662__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10475__A2 _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ _14472_/CLK _13878_/D vssd1 vssd1 vccd1 vccd1 _13878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10786__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _13394_/B _13104_/A2 _12828_/X vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13162__B _13162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12847__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10227__A2 _13397_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11424__A1 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B2 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_150_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _14791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _08091_/B _08020_/B _08020_/C vssd1 vssd1 vccd1 vccd1 _08095_/A sky130_fd_sc_hd__and3_1
XANTENNA__07587__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09368__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08272__A _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11188__B1 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold703 hold703/A vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 hold714/A vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold725 hold725/A vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 hold736/A vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 hold747/A vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 hold758/A vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _09971_/A _09971_/B vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold769 hold769/A vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07319__C _10951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13024__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__nand2_1
Xhold2104 _07046_/X vssd1 vssd1 vccd1 vccd1 _13862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2115 _13896_/Q vssd1 vssd1 vccd1 vccd1 hold2115/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2126 _07133_/X vssd1 vssd1 vccd1 vccd1 _13943_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12783__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2137 _14366_/Q vssd1 vssd1 vccd1 vccd1 hold2137/X sky130_fd_sc_hd__dlygate4sd3_1
X_08853_ _08744_/B _08746_/B _08742_/X vssd1 vssd1 vccd1 vccd1 _08854_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_209_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2148 _07087_/X vssd1 vssd1 vccd1 vccd1 _13900_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 _13986_/Q vssd1 vssd1 vccd1 vccd1 hold1403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 _11713_/X vssd1 vssd1 vccd1 vccd1 _14509_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2159 _14774_/Q vssd1 vssd1 vccd1 vccd1 hold2159/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08451__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1425 _13833_/Q vssd1 vssd1 vccd1 vccd1 hold1425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 _07202_/X vssd1 vssd1 vccd1 vccd1 _14009_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ hold547/X _11921_/A0 _07810_/S vssd1 vssd1 vccd1 vccd1 hold548/A sky130_fd_sc_hd__mux2_1
XANTENNA__11138__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1447 _14511_/Q vssd1 vssd1 vccd1 vccd1 hold1447/X sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ _09009_/A _09866_/B _08783_/C _08783_/D vssd1 vssd1 vccd1 vccd1 _08785_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13637__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1458 _07603_/X vssd1 vssd1 vccd1 vccd1 _14227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _15414_/Q vssd1 vssd1 vccd1 vccd1 hold1469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ hold1561/X _13741_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07735_/X sky130_fd_sc_hd__mux2_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13353__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ hold979/X _13705_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 hold980/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _10185_/A _09860_/B _09404_/C _09539_/A vssd1 vssd1 vccd1 vccd1 _09406_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout624_A _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07597_ hold103/X hold2818/X _07609_/S vssd1 vssd1 vccd1 vccd1 hold104/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _09762_/A _09762_/B _09202_/A vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09267_ _09724_/D _09124_/B _09127_/B vssd1 vssd1 vccd1 vccd1 _09269_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15384_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07497__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08218_ _08149_/A _08149_/C _08149_/B vssd1 vssd1 vccd1 vccd1 _08230_/A sky130_fd_sc_hd__o21bai_1
X_09198_ _09198_/A _09198_/B vssd1 vssd1 vccd1 vccd1 _09201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12376__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ _08149_/A _08149_/B _08149_/C vssd1 vssd1 vccd1 vccd1 _08152_/A sky130_fd_sc_hd__or3_1
XANTENNA__08044__B1 _14428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ _11160_/A _11160_/B _11160_/C vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__and3_1
XFILLER_0_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11747__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _10110_/A _14961_/Q _10280_/A _10110_/D vssd1 vssd1 vccd1 vccd1 _10111_/X
+ sky130_fd_sc_hd__a22o_1
X_11091_ _11091_/A _11091_/B vssd1 vssd1 vccd1 vccd1 _11093_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10042_ _10042_/A _10042_/B _10042_/C vssd1 vssd1 vccd1 vccd1 _10044_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12774__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09444__C _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11048__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2660 _14438_/Q vssd1 vssd1 vccd1 vccd1 _09087_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2671 _14817_/Q vssd1 vssd1 vccd1 vccd1 hold2671/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07245__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _15254_/CLK _14850_/D vssd1 vssd1 vccd1 vccd1 _14850_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2682 _14823_/Q vssd1 vssd1 vccd1 vccd1 hold2682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2693 _08543_/X vssd1 vssd1 vccd1 vccd1 _14434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ _15072_/CLK _13801_/D vssd1 vssd1 vccd1 vccd1 _13801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1970 _07013_/X vssd1 vssd1 vccd1 vccd1 _13830_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1981 _14459_/Q vssd1 vssd1 vccd1 vccd1 hold1981/X sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _15261_/CLK hold590/X vssd1 vssd1 vccd1 vccd1 hold589/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1992 _07616_/X vssd1 vssd1 vccd1 vccd1 _14239_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ hold369/X _13715_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 hold370/A sky130_fd_sc_hd__mux2_1
XFILLER_0_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13263__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_13732_ hold881/X _13732_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 hold882/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10457__A2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__B1 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ hold807/A _14553_/Q hold731/A _14777_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _10944_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13663_ hold1519/X _13663_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 _13663_/X sky130_fd_sc_hd__mux2_1
X_10875_ _10875_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10876_/B sky130_fd_sc_hd__and2_1
X_15402_ _15405_/CLK hold804/X vssd1 vssd1 vccd1 vccd1 hold803/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11406__A1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ hold611/X hold1933/X hold555/X hold1803/X _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12614_/X sky130_fd_sc_hd__mux4_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11406__B2 _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12603__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ _13594_/A _13636_/B vssd1 vssd1 vccd1 vccd1 _13594_/X sky130_fd_sc_hd__or2_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15333_ _15340_/CLK _15333_/D vssd1 vssd1 vccd1 vccd1 _15333_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11501__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ _12545_/A _12545_/B _12601_/A vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_132_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15451_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ _15264_/CLK _15264_/D vssd1 vssd1 vccd1 vccd1 _15264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12476_ _12676_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _12477_/C sky130_fd_sc_hd__or2_1
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07200__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12906__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ _14602_/CLK _14215_/D vssd1 vssd1 vccd1 vccd1 _14215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11427_ _11597_/A _14967_/Q _11427_/C _11574_/A vssd1 vssd1 vccd1 vccd1 _11574_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA_5 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15195_ _15384_/CLK _15195_/D vssd1 vssd1 vccd1 vccd1 _15195_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10917__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08130__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _14954_/CLK _14146_/D vssd1 vssd1 vccd1 vccd1 _14146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _11358_/A _11518_/B _11358_/C vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__and3_1
XANTENNA__12119__C1 _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ _10306_/Y _10307_/X _10131_/X _10134_/X vssd1 vssd1 vccd1 vccd1 _10310_/B
+ sky130_fd_sc_hd__a211o_1
X_14077_ _14077_/CLK _14077_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
X_11289_ _13749_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _11289_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13331__A1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__A1_N _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _13679_/A1 _12329_/B _13078_/B1 _13200_/B vssd1 vssd1 vccd1 vccd1 _13028_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13157__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10145__A1 _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10797__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14979_ _15250_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 _14979_/Q sky130_fd_sc_hd__dfxtp_1
X_07520_ hold1233/X _13691_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13173__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07451_ _07451_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _14081_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07382_ _13240_/A _14062_/Q _07405_/A _15350_/Q vssd1 vssd1 vccd1 vccd1 _07382_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _08841_/B _09117_/Y _09119_/Y _09120_/Y _09070_/Y vssd1 vssd1 vccd1 vccd1
+ _09762_/A sky130_fd_sc_hd__o2111a_2
XFILLER_0_146_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13070__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_123_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _14472_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _09049_/X _09050_/Y _08930_/B _08932_/B vssd1 vssd1 vccd1 vccd1 _09052_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07110__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08003_ hold2756/X input27/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13176_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold500 hold500/A vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 hold511/A vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold522 hold522/A vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold533 hold533/A vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold544 hold544/A vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 hold555/A vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 hold566/A vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold577 hold577/A vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 hold588/A vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13348__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09954_ _11320_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 hold599/A vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12252__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__A1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ _09816_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _08915_/A sky130_fd_sc_hd__nand2_1
X_09885_ _09888_/B vssd1 vssd1 vccd1 vccd1 _09885_/Y sky130_fd_sc_hd__inv_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout574_A _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1200 _07059_/X vssd1 vssd1 vccd1 vccd1 _13875_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 _14285_/Q vssd1 vssd1 vccd1 vccd1 hold1211/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08953_/A _08834_/X _08693_/Y _08696_/Y vssd1 vssd1 vccd1 vccd1 _08836_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 _13701_/X vssd1 vssd1 vccd1 vccd1 _15407_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 _14145_/Q vssd1 vssd1 vccd1 vccd1 hold1233/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1244 _11884_/X vssd1 vssd1 vccd1 vccd1 _14706_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07780__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1255 _15421_/Q vssd1 vssd1 vccd1 vccd1 hold1255/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09561__A _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1266 _07662_/X vssd1 vssd1 vccd1 vccd1 _14283_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12508__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _15403_/Q _14538_/Q _14698_/Q _14762_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08767_/X sky130_fd_sc_hd__mux4_1
Xhold1277 _13852_/Q vssd1 vssd1 vccd1 vccd1 hold1277/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13086__B1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1288 _07065_/X vssd1 vssd1 vccd1 vccd1 _13881_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1299 _13948_/Q vssd1 vssd1 vccd1 vccd1 hold1299/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout839_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08188__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ hold851/X _13724_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold852/A sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _08607_/A _08699_/B _08606_/B _08608_/B _08608_/A vssd1 vssd1 vccd1 vccd1
+ _08712_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07649_ hold1181/X _13721_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 _07649_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10660_ _10660_/A _10660_/B _10660_/C vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_193_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08905__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _09184_/B _09186_/B _09316_/Y _09318_/X vssd1 vssd1 vccd1 vccd1 _09321_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08265__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_114_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15410_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ _11497_/A _10591_/B vssd1 vssd1 vccd1 vccd1 _10591_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12427__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ _12330_/A _12330_/B vssd1 vssd1 vccd1 vccd1 _12330_/X sky130_fd_sc_hd__and2_4
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _13455_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _14910_/D sky130_fd_sc_hd__and2_1
XFILLER_0_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14000_ _15079_/CLK _14000_/D vssd1 vssd1 vccd1 vccd1 _14000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11212_ _11212_/A _11212_/B _11212_/C vssd1 vssd1 vccd1 vccd1 _11370_/A sky130_fd_sc_hd__and3_1
XFILLER_0_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12192_ _14907_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__or2_1
XANTENNA__08663__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _11578_/A _11577_/A _14968_/Q _14969_/Q vssd1 vssd1 vccd1 vccd1 _11146_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13313__A1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10127__A1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ _11070_/X _11071_/Y _10887_/X _10889_/Y vssd1 vssd1 vccd1 vccd1 _11076_/C
+ sky130_fd_sc_hd__a211oi_2
Xinput120 in1[30] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10127__B2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput131 in2[11] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13692__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput142 in2[21] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10025_ _10024_/B _10024_/C _10024_/A vssd1 vssd1 vccd1 vccd1 _10025_/Y sky130_fd_sc_hd__o21ai_1
X_14902_ _14987_/CLK _14902_/D vssd1 vssd1 vccd1 vccd1 _14902_/Q sky130_fd_sc_hd__dfxtp_1
Xinput153 in2[31] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__clkbuf_2
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07690__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2490 _12123_/X vssd1 vssd1 vccd1 vccd1 _14873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14833_ _14842_/CLK _14833_/D vssd1 vssd1 vccd1 vccd1 _14833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13616__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _15405_/CLK _14764_/D vssd1 vssd1 vccd1 vccd1 _14764_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ hold639/X _13665_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 hold640/A sky130_fd_sc_hd__mux2_1
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13715_ hold1255/X _13715_/A1 _13715_/S vssd1 vssd1 vccd1 vccd1 _13715_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11225__B _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ hold2357/X _07812_/A _13590_/B _10924_/Y _10926_/X vssd1 vssd1 vccd1 vccd1
+ _10927_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ _15437_/CLK hold430/X vssd1 vssd1 vccd1 vccd1 hold429/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11940__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13646_ input56/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13646_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10858_ _10673_/A _10673_/Y _11037_/B _10857_/X vssd1 vssd1 vccd1 vccd1 _10900_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12588__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_105_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _15247_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13577_ _09773_/B _13586_/B _13576_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13577_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10789_ _10790_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__and2b_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _15316_/CLK _15316_/D vssd1 vssd1 vccd1 vccd1 _15316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12528_ _13659_/A1 _12329_/B _12953_/B1 _13180_/B vssd1 vssd1 vccd1 vccd1 _12528_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _15247_/CLK hold90/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
X_12459_ hold1047/X hold2147/X _12459_/S vssd1 vssd1 vccd1 vccd1 _12459_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ _15371_/CLK _15178_/D vssd1 vssd1 vccd1 vccd1 _15178_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09220__A2 _12276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__D _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ _15196_/CLK _14129_/D vssd1 vssd1 vccd1 vccd1 _14129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13304__A1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12107__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _06950_/X _07453_/A _14029_/Q vssd1 vssd1 vccd1 vccd1 _06951_/X sky130_fd_sc_hd__and3b_4
XFILLER_0_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10304__B _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09670_ _10351_/A _10338_/C _09671_/A vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08621_ _08621_/A _08621_/B _08621_/C vssd1 vssd1 vccd1 vccd1 _08621_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13615__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08552_ _14792_/Q _14504_/Q _14632_/Q _14728_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08553_/B sky130_fd_sc_hd__mux4_1
XANTENNA__07105__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07503_ hold1475/X _11921_/A0 _07509_/S vssd1 vssd1 vccd1 vccd1 _07503_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08483_ _08483_/A _08483_/B _08483_/C vssd1 vssd1 vccd1 vccd1 _08581_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11850__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07434_ _08741_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14064_/D sky130_fd_sc_hd__and2_1
XFILLER_0_175_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10841__A2 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07365_ _15349_/Q _14062_/Q vssd1 vssd1 vccd1 vccd1 _07365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_162_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12247__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09104_ hold539/A hold545/A _14410_/Q _14122_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09105_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ _07296_/A _07296_/B vssd1 vssd1 vccd1 vccd1 _10951_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _09035_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07775__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__A1 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 hold341/A vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08460__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__B2 _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 hold352/A vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A _14941_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold363 hold363/A vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold374 hold374/A vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold385 hold385/A vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 hold396/A vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout810 _14489_/Q vssd1 vssd1 vccd1 vccd1 _12899_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout821 _14488_/Q vssd1 vssd1 vccd1 vccd1 _12460_/S sky130_fd_sc_hd__buf_6
Xfanout832 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _12791_/S sky130_fd_sc_hd__buf_6
X_09937_ _11497_/A _09936_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _09937_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10109__A1 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout843 _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__buf_4
XANTENNA__10109__B2 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _07448_/B vssd1 vssd1 vccd1 vccd1 _07450_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout865 _13479_/A vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__clkbuf_8
Xfanout876 _13479_/A vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__buf_4
X_09868_ _09715_/A _09715_/B _09715_/C vssd1 vssd1 vccd1 vccd1 _09869_/C sky130_fd_sc_hd__a21bo_1
Xfanout887 _13150_/A vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__buf_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _07019_/X vssd1 vssd1 vccd1 vccd1 _13836_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 _14704_/Q vssd1 vssd1 vccd1 vccd1 hold1041/X sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _08820_/A _08820_/B _08820_/C vssd1 vssd1 vccd1 vccd1 _08819_/X sky130_fd_sc_hd__and3_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _11904_/X vssd1 vssd1 vccd1 vccd1 _14725_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _13801_/Q vssd1 vssd1 vccd1 vccd1 hold1063/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ hold921/A _13947_/Q _15448_/Q _13915_/Q _10425_/S0 _10425_/S1 vssd1 vssd1
+ vccd1 vccd1 _09800_/B sky130_fd_sc_hd__mux4_1
Xhold1074 _07164_/X vssd1 vssd1 vccd1 vccd1 _13972_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _14801_/Q vssd1 vssd1 vccd1 vccd1 hold1085/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 _07739_/X vssd1 vssd1 vccd1 vccd1 _14358_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_203 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ hold2189/X _12329_/A _11845_/S vssd1 vssd1 vccd1 vccd1 _11830_/X sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12806__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_214 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__A2 _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07015__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _13714_/A1 hold1895/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11761_/X sky130_fd_sc_hd__mux2_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11760__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ _13501_/A hold113/X vssd1 vssd1 vccd1 vccd1 hold114/A sky130_fd_sc_hd__and2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10712_ _10709_/X _10710_/Y _10534_/X _10536_/Y vssd1 vssd1 vccd1 vccd1 _10713_/C
+ sky130_fd_sc_hd__a211oi_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _15408_/CLK _14480_/D vssd1 vssd1 vccd1 vccd1 _14480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _06904_/A _13792_/A2 _11691_/X _07475_/B vssd1 vssd1 vccd1 vccd1 _14491_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13431_ _08743_/A _13440_/S _13430_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15209_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ _11542_/A _11606_/A _11536_/A _10827_/C vssd1 vssd1 vccd1 vccd1 _10646_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_165_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10045__B1 _10044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13362_ _13369_/A _13362_/B vssd1 vssd1 vccd1 vccd1 _15153_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10574_ _13750_/A _13367_/B _10572_/X _10573_/Y vssd1 vssd1 vccd1 vccd1 _10574_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ _15116_/CLK _15101_/D vssd1 vssd1 vccd1 vccd1 _15101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13687__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ _14653_/Q _13926_/Q _15427_/Q _13894_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12313_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12591__S _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _13317_/A _13293_/B vssd1 vssd1 vccd1 vccd1 _15117_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07685__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ _15196_/CLK _15032_/D vssd1 vssd1 vccd1 vccd1 _15032_/Q sky130_fd_sc_hd__dfxtp_1
X_12244_ hold509/A hold497/A _14139_/Q _14457_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _12245_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12175_ hold2605/X _12195_/A2 _12174_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12175_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10405__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ _11497_/A _11123_/X _11125_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _11127_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11935__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__S1 _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _11541_/A _11351_/B _11564_/B _11614_/B _10881_/X vssd1 vssd1 vccd1 vccd1
+ _11065_/A sky130_fd_sc_hd__a41o_1
XANTENNA__11848__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ _15200_/Q _10115_/A _10283_/C _10115_/D vssd1 vssd1 vccd1 vccd1 _10010_/D
+ sky130_fd_sc_hd__nand4_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14816_ _14844_/CLK _14816_/D vssd1 vssd1 vccd1 vccd1 _14816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12766__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14747_ _15196_/CLK _14747_/D vssd1 vssd1 vccd1 vccd1 _14747_/Q sky130_fd_sc_hd__dfxtp_1
X_11959_ _13714_/A1 hold795/X _11959_/S vssd1 vssd1 vccd1 vccd1 hold796/A sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11670__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ _15415_/CLK _14678_/D vssd1 vssd1 vccd1 vccd1 _14678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13629_ hold2331/X _13797_/A2 _13628_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15342_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ _13651_/A1 hold2257/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07150_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _12329_/A hold1849/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07081_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07595__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10339__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08280__A _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10339__B2 _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07204__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11000__A2 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09526__D _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__A4 _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13289__B1 _13288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ hold185/A _14302_/Q hold861/A _13962_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07983_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_129_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06963__B1 _06959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11845__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _10002_/C _10010_/B _09562_/X _09427_/B _10115_/D vssd1 vssd1 vccd1 vccd1
+ _09729_/A sky130_fd_sc_hd__a32o_1
XANTENNA__13626__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ _14090_/Q vssd1 vssd1 vccd1 vccd1 _11729_/C sky130_fd_sc_hd__inv_2
XFILLER_0_198_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08704__A1 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09653_ hold2748/X input13/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13192_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09542__C _15209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08604_ _08926_/A _08702_/B _08604_/C _08699_/A vssd1 vssd1 vccd1 vccd1 _08699_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09584_ _10115_/B _09726_/B _09584_/C _09584_/D vssd1 vssd1 vccd1 vccd1 _09721_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_210_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08535_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08536_/B sky130_fd_sc_hd__or2_1
XANTENNA__10985__A _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout537_A _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13361__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08466_ hold2746/X input2/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13182_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07417_ hold11/X _07473_/B vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__and2_1
XFILLER_0_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08397_ _08397_/A _08397_/B _08397_/C vssd1 vssd1 vccd1 vccd1 _08468_/A sky130_fd_sc_hd__nand3_2
XANTENNA_fanout704_A _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _15355_/Q _15354_/Q _15353_/Q _15352_/Q vssd1 vssd1 vccd1 vccd1 _07351_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07279_ _15221_/Q _14965_/Q vssd1 vssd1 vccd1 vccd1 _07280_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09019_/B sky130_fd_sc_hd__nand2_1
X_10290_ _10114_/B _10120_/B _10114_/A vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10425__S1 _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout640 _15200_/Q vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__clkbuf_8
Xfanout651 _15197_/Q vssd1 vssd1 vccd1 vccd1 _08677_/A sky130_fd_sc_hd__buf_4
XANTENNA__11755__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 _13711_/A1 vssd1 vssd1 vccd1 vccd1 _13744_/A1 sky130_fd_sc_hd__clkbuf_4
X_13980_ _15063_/CLK _13980_/D vssd1 vssd1 vccd1 vccd1 _13980_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout673 _13739_/A1 vssd1 vssd1 vccd1 vccd1 _13673_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10879__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 _13734_/A1 vssd1 vssd1 vccd1 vccd1 _13668_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout695 _15049_/Q vssd1 vssd1 vccd1 vccd1 _13729_/A1 sky130_fd_sc_hd__buf_4
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _13106_/A1 _13164_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12932_/B sky130_fd_sc_hd__o21a_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__B _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _13074_/S1 _12859_/X _12861_/X vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__a21o_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ hold1383/X _13519_/A0 _11828_/S vssd1 vssd1 vccd1 vccd1 _11813_/X sky130_fd_sc_hd__mux2_1
X_14601_ _15432_/CLK _14601_/D vssd1 vssd1 vccd1 vccd1 _14601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11058__A2 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12255__A1 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12255__B2 _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ _12899_/S1 _12790_/X _12792_/X vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__a21o_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _15361_/CLK hold902/X vssd1 vssd1 vccd1 vccd1 hold901/A sky130_fd_sc_hd__dfxtp_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _13730_/A1 hold1501/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11744_/X sky130_fd_sc_hd__mux2_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07131__A0 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08365__A _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14463_ _15040_/CLK _14463_/D vssd1 vssd1 vccd1 vccd1 _14463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11675_ hold2819/X hold729/X _11684_/S vssd1 vssd1 vccd1 vccd1 hold730/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09959__B1 _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _13466_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _13414_/Y sky130_fd_sc_hd__nand2_1
X_10626_ _10623_/Y _10624_/X _10447_/X _10452_/A vssd1 vssd1 vccd1 vccd1 _10627_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_181_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ _15390_/CLK hold592/X vssd1 vssd1 vccd1 vccd1 hold591/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_output191_A _15172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12963__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13345_ _13369_/A _13345_/B vssd1 vssd1 vccd1 vccd1 _15136_/D sky130_fd_sc_hd__nor2_1
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13210__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ input131/X fanout6/X fanout4/X input99/X vssd1 vssd1 vccd1 vccd1 _13276_/X
+ sky130_fd_sc_hd__a22o_1
X_10488_ _11407_/A _11390_/A _10652_/A _10487_/D vssd1 vssd1 vccd1 vccd1 _10489_/C
+ sky130_fd_sc_hd__a22o_1
X_15015_ _15436_/CLK _15015_/D vssd1 vssd1 vccd1 vccd1 _15015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12227_ _13373_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _14909_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_209_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _14890_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12158_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11665__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ _10921_/B _10744_/B _11645_/A vssd1 vssd1 vccd1 vccd1 _11110_/B sky130_fd_sc_hd__o21a_1
X_12089_ hold2424/X _12099_/A2 _12088_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12089_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07444__A _08253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13165__B _13165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12494__A1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ _08320_/A _08320_/B _08413_/A _08320_/D vssd1 vssd1 vccd1 vccd1 _08322_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08251_ _08181_/A _08178_/Y _08180_/B vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07202_ hold1435/X _13703_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 _07202_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13746__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ hold2687/X _09925_/A2 _07390_/A vssd1 vssd1 vccd1 vccd1 _08182_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07133_ _13734_/A1 hold2125/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07133_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07064_ _13669_/A1 hold2091/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07064_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput210 _14192_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[22] sky130_fd_sc_hd__buf_12
XFILLER_0_30_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput221 _14173_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[3] sky130_fd_sc_hd__buf_12
Xoutput232 _14437_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[13] sky130_fd_sc_hd__buf_12
XFILLER_0_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput243 _14447_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[23] sky130_fd_sc_hd__buf_12
Xoutput254 _14428_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[4] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput265 _14891_/Q vssd1 vssd1 vccd1 vccd1 out0[14] sky130_fd_sc_hd__buf_12
Xoutput276 _14901_/Q vssd1 vssd1 vccd1 vccd1 out0[24] sky130_fd_sc_hd__buf_12
XFILLER_0_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput287 _14882_/Q vssd1 vssd1 vccd1 vccd1 out0[5] sky130_fd_sc_hd__buf_12
XFILLER_0_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput298 _14860_/Q vssd1 vssd1 vccd1 vccd1 out1[15] sky130_fd_sc_hd__buf_12
XFILLER_0_103_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13356__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _07965_/A _07964_/X _07965_/Y vssd1 vssd1 vccd1 vccd1 _07966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09705_ _09706_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09856_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_199_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06917_ hold261/X vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ hold2789/X _12256_/A _12258_/S _07896_/Y vssd1 vssd1 vccd1 vccd1 _07897_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _14975_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout654_A _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _10244_/A _09633_/X _09635_/X vssd1 vssd1 vccd1 vccd1 _09636_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09567_ _09708_/B _09430_/X _09566_/X vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_167_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout821_A _14488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08185__A _14430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _09498_/A _14442_/Q _09498_/C vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__and3_1
XFILLER_0_182_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ _12243_/A _08446_/X _08448_/X vssd1 vssd1 vccd1 vccd1 _08449_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11460_ _11460_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09405__A2 _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _15157_/Q _07812_/A _13634_/B _10410_/X vssd1 vssd1 vccd1 vccd1 _10411_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _11390_/A _11537_/B _11390_/C _11390_/D vssd1 vssd1 vccd1 vccd1 _11392_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ _13489_/A hold33/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__and2_1
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09169__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12399__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ _13092_/A1 _13060_/X _13100_/S0 vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07248__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10273_ _14964_/Q _10273_/B vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12012_ hold2653/X hold2667/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12013_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13266__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout470 _12128_/C vssd1 vssd1 vccd1 vccd1 _12096_/C sky130_fd_sc_hd__clkbuf_4
Xfanout492 _06944_/Y vssd1 vssd1 vccd1 vccd1 _12700_/S1 sky130_fd_sc_hd__buf_8
X_13963_ _15042_/CLK _13963_/D vssd1 vssd1 vccd1 vccd1 _13963_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_85_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _14926_/CLK sky130_fd_sc_hd__clkbuf_16
X_12914_ hold425/A _14226_/Q hold467/A _14480_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12914_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12571__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13894_ _15427_/CLK _13894_/D vssd1 vssd1 vccd1 vccd1 _13894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10582__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12845_ _12845_/A _12845_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__or3b_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13205__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12776_ _12951_/A _12776_/B vssd1 vssd1 vccd1 vccd1 _12777_/C sky130_fd_sc_hd__or2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07203__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12329__B _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11233__B _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ _15372_/CLK _14515_/D vssd1 vssd1 vccd1 vccd1 _14515_/Q sky130_fd_sc_hd__dfxtp_1
X_11727_ hold875/X _13681_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 hold876/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09919__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11658_ _13689_/A1 hold1141/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11658_/X sky130_fd_sc_hd__mux2_1
X_14446_ _15316_/CLK _14446_/D vssd1 vssd1 vccd1 vccd1 _14446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ _10609_/A _10788_/B vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__or2_1
XFILLER_0_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11203__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ _15373_/CLK _14377_/D vssd1 vssd1 vccd1 vccd1 _14377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11589_ _11598_/A _11573_/B _11441_/B vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold907 hold907/A vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ input85/X fanout2/X _13327_/X vssd1 vssd1 vccd1 vccd1 _13329_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10411__B1 _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold918 hold918/A vssd1 vssd1 vccd1 vccd1 hold918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold929 hold929/A vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10962__A1 _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ input92/X fanout1/X _13258_/X vssd1 vssd1 vccd1 vccd1 _13260_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12703__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2308 _14032_/Q vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2319 _14973_/Q vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09580__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13176__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _15360_/Q _15263_/Q _15071_/Q _14364_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _07820_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09580__B2 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2417_A _14070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1607 _15408_/Q vssd1 vssd1 vccd1 vccd1 hold1607/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1618 _11834_/X vssd1 vssd1 vccd1 vccd1 _14657_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1629 _14777_/Q vssd1 vssd1 vccd1 vccd1 hold1629/X sky130_fd_sc_hd__dlygate4sd3_1
X_07751_ _13656_/A1 hold2013/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07751_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12467__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15456_/CLK sky130_fd_sc_hd__clkbuf_16
X_07682_ hold1281/X _13655_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 _07682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09421_ _09421_/A vssd1 vssd1 vccd1 vccd1 _09421_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13623__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2786_A _15195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11690__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12314__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _10233_/A _09498_/C _09352_/C vssd1 vssd1 vccd1 vccd1 _09352_/X sky130_fd_sc_hd__or3_1
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ _09661_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__and2_1
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11143__B _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_150_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09283_ _10338_/B _09860_/B _09676_/D _10166_/A vssd1 vssd1 vccd1 vccd1 _09285_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _08234_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_30_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10982__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ _08240_/A _08164_/C _08164_/A vssd1 vssd1 vccd1 vccd1 _08165_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_16_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout402_A _07477_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10402__B1 _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_165_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07116_ _12329_/A hold2285/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07116_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08071__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08096_ _08095_/B _08095_/C _08095_/A vssd1 vssd1 vccd1 vccd1 _08097_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_45_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ _13652_/A1 hold1653/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07047_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07783__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2820 _15340_/Q vssd1 vssd1 vccd1 vccd1 hold2820/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2831 _15318_/Q vssd1 vssd1 vccd1 vccd1 hold2831/X sky130_fd_sc_hd__dlygate4sd3_1
X_08998_ _09846_/B _09726_/B _09724_/C _10000_/A vssd1 vssd1 vccd1 vccd1 _09001_/A
+ sky130_fd_sc_hd__a22o_1
Xhold2842 _15332_/Q vssd1 vssd1 vccd1 vccd1 hold2842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2853 _15310_/Q vssd1 vssd1 vccd1 vccd1 hold2853/X sky130_fd_sc_hd__dlygate4sd3_1
X_07949_ _13687_/A1 _12260_/A2 _12259_/A1 _13175_/B _07947_/Y vssd1 vssd1 vccd1 vccd1
+ _07949_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14042_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10469__B1 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_103_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _10734_/A _10910_/X _10958_/X _10735_/Y _10912_/B vssd1 vssd1 vccd1 vccd1
+ _10960_/X sky130_fd_sc_hd__o221a_2
XFILLER_0_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08908__A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09874__A2 _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07812__A _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ _09619_/A _09619_/B _09619_/C vssd1 vssd1 vccd1 vccd1 _09619_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_211_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10891_ _10707_/Y _10709_/X _10889_/Y _10890_/X vssd1 vssd1 vccd1 vccd1 _10893_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ _12327_/A _12629_/X _12627_/X vssd1 vssd1 vccd1 vccd1 _13152_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__B _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ _12692_/A1 _12560_/X _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12630__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14300_ _15263_/CLK hold302/X vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
X_11512_ _12252_/B _11512_/B vssd1 vssd1 vccd1 vccd1 _11512_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15280_ _15377_/CLK _15280_/D vssd1 vssd1 vccd1 vccd1 _15280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12492_ _12642_/A1 _12491_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _15456_/CLK _14231_/D vssd1 vssd1 vccd1 vccd1 _14231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11443_ _11443_/A _11443_/B _11443_/C vssd1 vssd1 vccd1 vccd1 _11445_/C sky130_fd_sc_hd__and3_1
XFILLER_0_180_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07259__A _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _15451_/CLK hold468/X vssd1 vssd1 vccd1 vccd1 hold467/A sky130_fd_sc_hd__dfxtp_1
X_11374_ _11374_/A _11374_/B vssd1 vssd1 vccd1 vccd1 _11376_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13695__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ _13129_/A hold45/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__and2_1
X_10325_ _10324_/A _10324_/B _10324_/C vssd1 vssd1 vccd1 vccd1 _10326_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14093_ _14105_/CLK hold274/X vssd1 vssd1 vccd1 vccd1 _14093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09237__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13100_/S0 _13039_/X _13043_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _13045_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _10241_/Y _10246_/Y _10255_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _10257_/B sky130_fd_sc_hd__a221o_1
XANTENNA__09562__A1 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09562__B2 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _10019_/D _10020_/B _10185_/X _10186_/Y vssd1 vssd1 vccd1 vccd1 _10189_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08770__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15127_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10132__B _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14995_ _15248_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 _14995_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11943__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ _15448_/CLK _13946_/D vssd1 vssd1 vccd1 vccd1 _13946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11121__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07876__A1 _15341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _14409_/CLK _13877_/D vssd1 vssd1 vccd1 vccd1 _13877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10880__B1 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _13704_/A1 _13103_/A2 _13078_/B1 _13192_/B vssd1 vssd1 vccd1 vccd1 _12828_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11424__A2 _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ hold427/A _13912_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08553__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14429_ _15299_/CLK _14429_/D vssd1 vssd1 vccd1 vccd1 _14429_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11188__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08053__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold704 hold704/A vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold715 hold715/A vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 hold726/A vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 hold737/A vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _09971_/A _09971_/B vssd1 vssd1 vccd1 vccd1 _09970_/Y sky130_fd_sc_hd__nand2_1
Xhold748 hold748/A vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 hold759/A vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07319__D _07319_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09384__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ _08788_/A _08787_/B _08785_/X vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12688__A1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2105 _14140_/Q vssd1 vssd1 vccd1 vccd1 hold2105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2701_A _14843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2116 _07083_/X vssd1 vssd1 vccd1 vccd1 _13896_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10699__B1 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2127 _14760_/Q vssd1 vssd1 vccd1 vccd1 hold2127/X sky130_fd_sc_hd__dlygate4sd3_1
X_08852_ _08850_/X _08852_/B vssd1 vssd1 vccd1 vccd1 _08854_/A sky130_fd_sc_hd__and2b_1
Xhold2138 _07750_/X vssd1 vssd1 vccd1 vccd1 _14366_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12783__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1404 _07178_/X vssd1 vssd1 vccd1 vccd1 _13986_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2149 _15271_/Q vssd1 vssd1 vccd1 vccd1 hold2149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 _14410_/Q vssd1 vssd1 vccd1 vccd1 hold1415/X sky130_fd_sc_hd__dlygate4sd3_1
X_07803_ hold897/X _13741_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold898/A sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07108__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1426 _07016_/X vssd1 vssd1 vccd1 vccd1 _13833_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ _09009_/A _09866_/B _08783_/C _08783_/D vssd1 vssd1 vccd1 vccd1 _08785_/B
+ sky130_fd_sc_hd__nand4_1
Xhold1437 _14604_/Q vssd1 vssd1 vccd1 vccd1 hold1437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1448 _11715_/X vssd1 vssd1 vccd1 vccd1 _14511_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15424_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1459 _13965_/Q vssd1 vssd1 vccd1 vccd1 hold1459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11853__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07734_ hold1369/X _13740_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07734_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07665_ hold805/X _13737_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 hold806/A sky130_fd_sc_hd__mux2_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _10185_/A _09860_/B _09404_/C _09539_/A vssd1 vssd1 vccd1 vccd1 _09539_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ _15055_/Q hold1905/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07596_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09762_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12612__A1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12684__S _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A _15205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09266_ _09449_/B _09266_/B vssd1 vssd1 vccd1 vccd1 _09269_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08217_ _08301_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__or2_1
XFILLER_0_132_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ _09198_/A _09198_/B vssd1 vssd1 vccd1 vccd1 _09197_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08148_ _08147_/A _08147_/B _08147_/C vssd1 vssd1 vccd1 vccd1 _08149_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__08044__A1 _14427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12471__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08007_/A _08007_/C _08007_/B vssd1 vssd1 vccd1 vccd1 _08080_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09294__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _10110_/A _14961_/Q _10280_/A _10110_/D vssd1 vssd1 vccd1 vccd1 _10280_/B
+ sky130_fd_sc_hd__nand4_2
X_11090_ _11273_/B _11090_/B vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12679__A1 _13388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09544__A1 _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _10042_/A _10042_/B _10042_/C vssd1 vssd1 vccd1 vccd1 _10041_/X sky130_fd_sc_hd__and3_1
XANTENNA__12774__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__A _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09444__D _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07018__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2650 _09356_/X vssd1 vssd1 vccd1 vccd1 _14441_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11048__B _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2661 _08974_/X vssd1 vssd1 vccd1 vccd1 _14438_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2672 _14825_/Q vssd1 vssd1 vccd1 vccd1 hold2672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2683 _12020_/X vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2694 _15167_/Q vssd1 vssd1 vccd1 vccd1 hold2694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1960 _11660_/X vssd1 vssd1 vccd1 vccd1 _14463_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13544__A _14428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _14783_/CLK _13800_/D vssd1 vssd1 vccd1 vccd1 _13800_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11639__C1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1971 _14003_/Q vssd1 vssd1 vccd1 vccd1 hold1971/X sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ hold2237/X _13681_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11992_/X sky130_fd_sc_hd__mux2_1
X_14780_ _15455_/CLK _14780_/D vssd1 vssd1 vccd1 vccd1 _14780_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11103__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1982 _11656_/X vssd1 vssd1 vccd1 vccd1 _14459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1993 _14723_/Q vssd1 vssd1 vccd1 vccd1 hold1993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10943_ _11504_/A _10943_/B vssd1 vssd1 vccd1 vccd1 _10943_/Y sky130_fd_sc_hd__nor2_1
X_13731_ hold1395/X hold2801/X _13732_/S vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10874_ _10875_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10876_/A sky130_fd_sc_hd__nor2_1
X_13662_ hold471/X _13662_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold472/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15438_/CLK hold778/X vssd1 vssd1 vccd1 vccd1 hold777/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ _12642_/B1 _12608_/X _12612_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12620_/A
+ sky130_fd_sc_hd__o211a_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11406__A2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13593_ _11106_/B _11650_/B _13592_/X _13459_/A vssd1 vssd1 vccd1 vccd1 _13593_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07688__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15332_ _15340_/CLK _15332_/D vssd1 vssd1 vccd1 vccd1 _15332_/Q sky130_fd_sc_hd__dfxtp_1
X_12544_ _06943_/Y _12539_/X _12543_/X _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12545_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08283__A1 _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12475_ _12471_/X _12472_/X _12474_/X _12473_/X _12644_/A1 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12476_/B sky130_fd_sc_hd__mux4_1
X_15263_ _15263_/CLK _15263_/D vssd1 vssd1 vccd1 vccd1 _15263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10408__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11426_ _11597_/A _14967_/Q _11427_/C _11574_/A vssd1 vssd1 vccd1 vccd1 _11431_/A
+ sky130_fd_sc_hd__a22o_1
X_14214_ _14731_/CLK _14214_/D vssd1 vssd1 vccd1 vccd1 _14214_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12906__A2 _13163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _15289_/CLK _15194_/D vssd1 vssd1 vccd1 vccd1 _15194_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output271_A _14878_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__A1 _10951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14145_ _15040_/CLK _14145_/D vssd1 vssd1 vccd1 vccd1 _14145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08130__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09783__A1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11938__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ _11518_/A _11356_/C _11356_/A vssd1 vssd1 vccd1 vccd1 _11358_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _10131_/X _10134_/X _10306_/Y _10307_/X vssd1 vssd1 vccd1 vccd1 _10308_/X
+ sky130_fd_sc_hd__o211a_1
X_14076_ _15356_/CLK _14076_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13438__B _13438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11288_ _11288_/A1 _13403_/B _11140_/X vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__a21oi_4
X_13027_ _13027_/A _13027_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__and3_1
X_10239_ _13886_/Q _14014_/Q _13854_/Q _13822_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10239_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11673__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09299__B1 _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ _15250_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 _14978_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10797__B _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13173__B _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12842__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ _15434_/CLK _13929_/D vssd1 vssd1 vccd1 vccd1 _13929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07450_ hold77/X _07450_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__and2_1
XFILLER_0_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07381_ _14051_/Q _07846_/A _07381_/C _07381_/D vssd1 vssd1 vccd1 vccd1 _07879_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_0_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ _09071_/A _09071_/B _08954_/X vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07598__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10605__B1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _08930_/B _08932_/B _09049_/X _09050_/Y vssd1 vssd1 vccd1 vccd1 _09051_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_155_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12358__B1 _13141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08002_ _12252_/B _08002_/B vssd1 vssd1 vccd1 vccd1 _08002_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold501 hold501/A vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold512 hold512/A vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 hold523/A vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold534 hold534/A vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09826__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 hold545/A vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold556 hold556/A vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08982__C1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 hold567/A vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 hold578/A vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _09938_/Y _09943_/Y _09952_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09954_/B sky130_fd_sc_hd__a221o_1
Xhold589 hold589/A vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12252__B _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ _08800_/A _08799_/B _08799_/A vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__o21ba_1
X_09884_ _09886_/A _09886_/B _09886_/C vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10136__A2 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _14456_/Q vssd1 vssd1 vccd1 vccd1 hold1201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _07664_/X vssd1 vssd1 vccd1 vccd1 _14285_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08835_ _08693_/Y _08696_/Y _08953_/A _08834_/X vssd1 vssd1 vccd1 vccd1 _08953_/B
+ sky130_fd_sc_hd__a211oi_2
Xhold1223 _14466_/Q vssd1 vssd1 vccd1 vccd1 hold1223/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1234 _07520_/X vssd1 vssd1 vccd1 vccd1 _14145_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout567_A _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 _14615_/Q vssd1 vssd1 vccd1 vccd1 hold1245/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13364__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 _13715_/X vssd1 vssd1 vccd1 vccd1 _15421_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09561__B _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08989_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08766_/Y sky130_fd_sc_hd__nor2_1
Xhold1267 _14709_/Q vssd1 vssd1 vccd1 vccd1 hold1267/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13086__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1278 _07035_/X vssd1 vssd1 vccd1 vccd1 _13852_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08458__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1289 _14691_/Q vssd1 vssd1 vccd1 vccd1 hold1289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08188__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ hold337/X _13690_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold338/A sky130_fd_sc_hd__mux2_1
X_08697_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _08717_/A sky130_fd_sc_hd__xnor2_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout734_A _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07648_ hold423/X _13687_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold424/A sky130_fd_sc_hd__mux2_1
XFILLER_0_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07579_ _13718_/A1 hold497/X _07593_/S vssd1 vssd1 vccd1 vccd1 hold498/A sky130_fd_sc_hd__mux2_1
XANTENNA__08905__B _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09318_ _09317_/B _09317_/C _09317_/A vssd1 vssd1 vccd1 vccd1 _09318_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_192_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08193__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10590_ _14679_/Q _13952_/Q hold833/A _13920_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _10591_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_146_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09249_ _10126_/A _09248_/X _09247_/X vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08360__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10228__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12349__B1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _13718_/A1 _12260_/A2 _12252_/Y _12259_/X vssd1 vssd1 vccd1 vccd1 _12261_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ _11022_/A _11022_/C _11022_/B vssd1 vssd1 vccd1 vccd1 _11212_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11758__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12191_ hold2542/X _12195_/A2 _12190_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12191_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11142_ _11577_/A _14968_/Q _14969_/Q _11578_/A vssd1 vssd1 vccd1 vccd1 _11146_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09517__A1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11076_/B vssd1 vssd1 vccd1 vccd1 _11073_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12747__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput110 in1[21] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10127__A2 _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput121 in1[31] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10758__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput132 in2[12] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__clkbuf_2
X_10024_ _10024_/A _10024_/B _10024_/C vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__or3_1
X_14901_ _14987_/CLK _14901_/D vssd1 vssd1 vccd1 vccd1 _14901_/Q sky130_fd_sc_hd__dfxtp_1
Xinput143 in2[22] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__clkbuf_2
Xinput154 in2[3] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__clkbuf_2
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2480 _14433_/Q vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__buf_1
XFILLER_0_192_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _14840_/CLK _14832_/D vssd1 vssd1 vccd1 vccd1 _14832_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2491 _14872_/Q vssd1 vssd1 vccd1 vccd1 hold2491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07272__A _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1790 _07062_/X vssd1 vssd1 vccd1 vccd1 _13878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _15367_/CLK _14763_/D vssd1 vssd1 vccd1 vccd1 _14763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ hold785/X _13664_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 hold786/A sky130_fd_sc_hd__mux2_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ hold783/X _13714_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold784/A sky130_fd_sc_hd__mux2_1
XFILLER_0_196_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11225__C _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10926_ _14451_/Q _11113_/C _10925_/Y _07390_/A vssd1 vssd1 vccd1 vccd1 _10926_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14694_ _15045_/CLK hold580/X vssd1 vssd1 vccd1 vccd1 hold579/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10930__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13645_ _08435_/A _13792_/A2 _13644_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15355_/D
+ sky130_fd_sc_hd__o211a_1
X_10857_ _11037_/A _10856_/B _10856_/C _10856_/D vssd1 vssd1 vccd1 vccd1 _10857_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13213__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10788_/A _10788_/B vssd1 vssd1 vccd1 vccd1 _10790_/B sky130_fd_sc_hd__or2_1
XFILLER_0_27_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _14444_/Q _13590_/B vssd1 vssd1 vccd1 vccd1 _13576_/X sky130_fd_sc_hd__or2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12683__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07211__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15315_ _15315_/CLK _15315_/D vssd1 vssd1 vccd1 vccd1 _15315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12527_ _13027_/A _12527_/B _12527_/C vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__and3_1
XFILLER_0_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09927__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15246_ _15246_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12458_ hold641/X hold2007/X _14691_/Q hold1445/X _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12458_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11668__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ _11409_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11410_/B sky130_fd_sc_hd__nand2_1
X_12389_ hold423/A _14205_/Q hold359/A _14459_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux4_1
X_15177_ _15177_/CLK _15177_/D vssd1 vssd1 vccd1 vccd1 _15177_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07447__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ _15062_/CLK _14128_/D vssd1 vssd1 vccd1 vccd1 _14128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06950_ _14030_/Q _06950_/B _06950_/C vssd1 vssd1 vccd1 vccd1 _06950_/X sky130_fd_sc_hd__or3_1
X_14059_ _15348_/CLK _14059_/D vssd1 vssd1 vccd1 vccd1 _14059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ _08617_/Y _08618_/X _08508_/Y _08510_/Y vssd1 vssd1 vccd1 vccd1 _08621_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13184__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08278__A _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09367__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ hold471/A hold705/A hold981/A _14373_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08551_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07502_ hold1683/X _13741_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07502_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08482_ _08389_/A _08389_/C _08389_/B vssd1 vssd1 vccd1 vccd1 _08483_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07433_ _07433_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _14063_/D sky130_fd_sc_hd__and2_1
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08247__A1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07364_ _15350_/Q _14063_/Q vssd1 vssd1 vccd1 vccd1 _07364_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_190_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12674__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09103_ _10246_/A _09103_/B vssd1 vssd1 vccd1 vccd1 _09103_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07121__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07295_ _15223_/Q _07295_/B vssd1 vssd1 vccd1 vccd1 _07296_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13791__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09034_ _09035_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _09034_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13359__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12263__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A2 _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 hold342/A vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/A vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 hold364/A vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold375/A vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout800 _12689_/S1 vssd1 vssd1 vccd1 vccd1 _12599_/S1 sky130_fd_sc_hd__clkbuf_8
Xhold386 hold386/A vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 hold397/A vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _12939_/S1 vssd1 vssd1 vccd1 vccd1 _06942_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout822 _12641_/S vssd1 vssd1 vccd1 vccd1 _12591_/S sky130_fd_sc_hd__buf_8
X_09936_ _13884_/Q hold675/A _13852_/Q _13820_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _09936_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout833 _12915_/S vssd1 vssd1 vccd1 vccd1 _12841_/S sky130_fd_sc_hd__buf_6
Xfanout844 _13565_/C1 vssd1 vssd1 vccd1 vccd1 _13579_/C1 sky130_fd_sc_hd__buf_4
Xfanout855 _13622_/C1 vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout866 _13490_/A vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__buf_4
Xfanout877 _12063_/A vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__buf_2
X_09867_ _10022_/B _09866_/B _09866_/C _09866_/D vssd1 vssd1 vccd1 vccd1 _09869_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout851_A _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout888 _13390_/A vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__clkbuf_8
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _07009_/X vssd1 vssd1 vccd1 vccd1 _13828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 _15079_/Q vssd1 vssd1 vccd1 vccd1 hold1031/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 _11882_/X vssd1 vssd1 vccd1 vccd1 _14704_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _08816_/B _08816_/C _08816_/A vssd1 vssd1 vccd1 vccd1 _08820_/C sky130_fd_sc_hd__a21o_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 _14787_/Q vssd1 vssd1 vccd1 vccd1 hold1053/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 _06982_/X vssd1 vssd1 vccd1 vccd1 _13801_/D sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _10426_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09798_/Y sky130_fd_sc_hd__nor2_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07930__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1075 _14920_/Q vssd1 vssd1 vccd1 vccd1 _13481_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09358__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1086 _11982_/X vssd1 vssd1 vccd1 vccd1 _14801_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1097 _15073_/Q vssd1 vssd1 vccd1 vccd1 hold1097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12806__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _09494_/A1 _08647_/Y _08748_/X vssd1 vssd1 vccd1 vccd1 _08749_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _13746_/A1 hold2199/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11760_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10711_ _10534_/X _10536_/Y _10709_/X _10710_/Y vssd1 vssd1 vccd1 vccd1 _10713_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__B1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11691_ input48/X _13648_/B vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__or2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10642_ _11542_/A _11606_/A _14954_/Q _10827_/C vssd1 vssd1 vccd1 vccd1 _10642_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_119_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13430_ _13440_/S _13430_/B vssd1 vssd1 vccd1 vccd1 _13430_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_193_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07031__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13361_ _13369_/A _13361_/B vssd1 vssd1 vccd1 vccd1 _15152_/D sky130_fd_sc_hd__nor2_1
X_10573_ _15158_/Q _07812_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _10573_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11793__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15100_ _15292_/CLK hold536/X vssd1 vssd1 vccd1 vccd1 hold535/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12312_ hold619/A _14202_/Q hold391/A _14456_/Q _12365_/S0 _12343_/A vssd1 vssd1
+ vccd1 vccd1 _12312_/X sky130_fd_sc_hd__mux4_1
X_13292_ input72/X fanout2/X _13291_/X vssd1 vssd1 vccd1 vccd1 _13293_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13269__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10108__D _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ _15063_/CLK _15031_/D vssd1 vssd1 vccd1 vccd1 _15031_/Q sky130_fd_sc_hd__dfxtp_1
X_12243_ _12243_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12742__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12174_ _14898_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__or2_1
XANTENNA__10405__B _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10753__C1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ _11507_/A _11125_/B vssd1 vssd1 vccd1 vccd1 _11125_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13298__A1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12901__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ _10835_/A _10834_/B _10832_/X vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__a21o_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _10110_/A _10115_/A _10283_/C _10115_/D vssd1 vssd1 vccd1 vccd1 _10007_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__13208__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11517__A _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07206__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _14876_/CLK _14815_/D vssd1 vssd1 vccd1 vccd1 _14815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11951__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14746_ _15387_/CLK _14746_/D vssd1 vssd1 vccd1 vccd1 _14746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11958_ _13746_/A1 hold1217/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__A1 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ _11098_/A _10907_/X _10690_/X _10693_/Y vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10284__B2 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14677_ _15093_/CLK hold772/X vssd1 vssd1 vccd1 vccd1 hold771/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11889_ hold1533/X _13743_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_157_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08229__A1 _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ input40/X _13634_/B vssd1 vssd1 vccd1 vccd1 _13628_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09977__A1 _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09977__B2 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ _08640_/A _09222_/B _13558_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _15305_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__B1 _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ _11652_/A _07115_/A vssd1 vssd1 vccd1 vccd1 _07080_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_129_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08561__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15229_ _15229_/CLK hold246/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13179__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10339__A2 _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07982_ _08042_/B _13591_/A2 _07970_/Y _07981_/X _13541_/A vssd1 vssd1 vccd1 vccd1
+ _07982_/X sky130_fd_sc_hd__o221a_1
X_09721_ _09721_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__nor2_1
X_06933_ _14089_/Q vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__inv_2
XFILLER_0_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13626__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08704__A2 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__A _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _11320_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09652_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09542__D _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07116__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _08776_/B _09138_/A _08809_/B _08809_/D vssd1 vssd1 vccd1 vccd1 _08699_/A
+ sky130_fd_sc_hd__nand4_2
X_09583_ _10115_/B _09726_/B _09584_/C _09584_/D vssd1 vssd1 vccd1 vccd1 _09585_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_96_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11861__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13642__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08534_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10985__B _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ _12252_/B _08465_/B vssd1 vssd1 vccd1 vccd1 _08465_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout432_A _11763_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07416_ hold15/X _07473_/B vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__and2_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08396_ _09816_/A _08685_/C _08395_/C _08395_/D vssd1 vssd1 vccd1 vccd1 _08397_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12647__S0 _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__B1 _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ _07362_/B _07362_/C vssd1 vssd1 vccd1 vccd1 _07351_/A sky130_fd_sc_hd__or2_1
XANTENNA__07786__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07278_ _15221_/Q _14965_/Q vssd1 vssd1 vccd1 vccd1 _07280_/A sky130_fd_sc_hd__or2_1
XFILLER_0_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09017_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__or2_1
XFILLER_0_143_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13072__S0 _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__buf_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout630 _15202_/Q vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__clkbuf_8
Xfanout641 _08075_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__buf_4
XANTENNA__07815__A _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout652 _15197_/Q vssd1 vssd1 vccd1 vccd1 _11580_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13536__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _10744_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09929_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12488__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout663 _15064_/Q vssd1 vssd1 vccd1 vccd1 _13711_/A1 sky130_fd_sc_hd__buf_4
Xfanout674 _15059_/Q vssd1 vssd1 vccd1 vccd1 _13739_/A1 sky130_fd_sc_hd__buf_4
Xfanout685 hold169/X vssd1 vssd1 vccd1 vccd1 _13734_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__10879__C _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout696 _13662_/A1 vssd1 vssd1 vccd1 vccd1 _13728_/A1 sky130_fd_sc_hd__clkbuf_4
X_12930_ _13080_/A1 _12929_/X _12927_/X vssd1 vssd1 vccd1 vccd1 _13164_/B sky130_fd_sc_hd__a21oi_4
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07026__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ _12917_/A1 _12860_/X _13100_/S0 vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__a21o_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11771__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12920__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _15268_/CLK _14600_/D vssd1 vssd1 vccd1 vccd1 _14600_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13552__A _14432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ hold1685/X _13666_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__mux2_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12255__A2 _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12792_ _12917_/A1 _12791_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__a21o_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07550__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14531_ _15433_/CLK _14531_/D vssd1 vssd1 vccd1 vccd1 _14531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _13729_/A1 hold2265/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11743_/X sky130_fd_sc_hd__mux2_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _15364_/CLK _14462_/D vssd1 vssd1 vccd1 vccd1 _14462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11674_ _13705_/A1 hold1777/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10018__A1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13698__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09959__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ _07974_/A _13450_/A _13412_/Y _13178_/A vssd1 vssd1 vccd1 vccd1 _15200_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09959__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10625_ _10447_/X _10452_/A _10623_/Y _10624_/X vssd1 vssd1 vccd1 vccd1 _10795_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14393_ _15292_/CLK _14393_/D vssd1 vssd1 vccd1 vccd1 _14393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07696__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11310__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10556_ _10553_/X _10554_/Y _10382_/Y _10387_/A vssd1 vssd1 vccd1 vccd1 _10557_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13344_ _13369_/A _13344_/B vssd1 vssd1 vccd1 vccd1 _15135_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output184_A _15167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ _13287_/A _13275_/B vssd1 vssd1 vccd1 vccd1 _15111_/D sky130_fd_sc_hd__nor2_1
X_10487_ _11407_/A _11390_/A _10652_/A _10487_/D vssd1 vssd1 vccd1 vccd1 _10652_/B
+ sky130_fd_sc_hd__nand4_2
X_15014_ _15177_/CLK _15014_/D vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__dfxtp_1
X_12226_ _12329_/A _12260_/A2 _12225_/X vssd1 vssd1 vccd1 vccd1 _13749_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__10135__B _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__A1 hold2542/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11946__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _14985_/Q _12173_/A2 _12156_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10741__A2 _11474_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _11108_/A _11108_/B _11108_/C _11108_/D vssd1 vssd1 vccd1 vccd1 _11111_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13446__B _13446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12088_ _14984_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12088_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__11247__A _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ _11081_/A vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07444__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13691__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11681__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13181__B _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ _15440_/CLK _14729_/D vssd1 vssd1 vccd1 vccd1 _14729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12078__A _14979_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08250_ _09918_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_184_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08870__A1 _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07201_ hold1055/X _13669_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 _07201_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _13348_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_hold2564_A _15001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11301__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ _13700_/A1 hold2183/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07132_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08291__A _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07063_ _13668_/A1 hold1723/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07063_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10326__A _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput200 _14183_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[13] sky130_fd_sc_hd__buf_12
Xoutput211 _14193_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[23] sky130_fd_sc_hd__buf_12
XFILLER_0_140_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12706__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput222 _14174_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[4] sky130_fd_sc_hd__buf_12
Xoutput233 _14438_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[14] sky130_fd_sc_hd__buf_12
XFILLER_0_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput244 _14448_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[24] sky130_fd_sc_hd__buf_12
XFILLER_0_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput255 _14429_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[5] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput266 _14892_/Q vssd1 vssd1 vccd1 vccd1 out0[15] sky130_fd_sc_hd__buf_12
XANTENNA__11856__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput277 _14902_/Q vssd1 vssd1 vccd1 vccd1 out0[25] sky130_fd_sc_hd__buf_12
Xoutput288 _14883_/Q vssd1 vssd1 vccd1 vccd1 out0[6] sky130_fd_sc_hd__buf_12
Xoutput299 _14861_/Q vssd1 vssd1 vccd1 vccd1 out1[16] sky130_fd_sc_hd__buf_12
XFILLER_0_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07965_ _07965_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _07965_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout382_A _11960_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09704_ _09704_/A _09704_/B vssd1 vssd1 vccd1 vccd1 _09706_/B sky130_fd_sc_hd__nor2_1
X_06916_ _06916_/A vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__inv_2
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ _07893_/Y _07895_/A _12256_/A vssd1 vssd1 vccd1 vccd1 _07896_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13682__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__A _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09635_ _10426_/A _09634_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _09635_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A1 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout647_A _15198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13372__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ _10126_/A _09708_/B _10126_/B _10022_/A vssd1 vssd1 vccd1 vccd1 _09566_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08517_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09497_ _14442_/Q _09498_/C _09498_/A vssd1 vssd1 vccd1 vccd1 _09497_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout814_A _14489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08185__B _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08448_ _12247_/A _08447_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08448_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08379_ _08378_/A _08378_/B _12258_/S vssd1 vssd1 vccd1 vccd1 _08379_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _13584_/A _10409_/B _10571_/B _07390_/A vssd1 vssd1 vccd1 vccd1 _10410_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11390_ _11390_/A _11537_/B _11390_/C _11390_/D vssd1 vssd1 vccd1 vccd1 _11392_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _11335_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09169__A2 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ hold487/A _13956_/Q _13066_/S vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__mux2_1
X_10272_ _11594_/B _10273_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12011_ _12063_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _14818_/D sky130_fd_sc_hd__and2_1
XANTENNA__12173__A1 hold2591/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10184__B1 _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07545__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout460 _12178_/B vssd1 vssd1 vccd1 vccd1 _12194_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout471 _12128_/C vssd1 vssd1 vccd1 vccd1 _12126_/C sky130_fd_sc_hd__clkbuf_4
Xfanout482 _07862_/X vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__buf_8
X_13962_ _14595_/CLK _13962_/D vssd1 vssd1 vccd1 vccd1 _13962_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout493 _13100_/S1 vssd1 vssd1 vccd1 vccd1 _12944_/C1 sky130_fd_sc_hd__buf_8
XANTENNA__11684__A0 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _12917_/B1 _12908_/X _12912_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12920_/A
+ sky130_fd_sc_hd__o211a_1
X_13893_ _15387_/CLK _13893_/D vssd1 vssd1 vccd1 vccd1 _13893_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10582__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12844_ _12844_/A1 _12839_/X _12843_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12845_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09629__B1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12775_ _12771_/X _12772_/X _12774_/X _12773_/X _12844_/A1 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12776_/B sky130_fd_sc_hd__mux4_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11987__A1 _15062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14514_ _15379_/CLK _14514_/D vssd1 vssd1 vccd1 vccd1 _14514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11726_ hold413/X _13680_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 hold414/A sky130_fd_sc_hd__mux2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14445_ _15315_/CLK _14445_/D vssd1 vssd1 vccd1 vccd1 _14445_/Q sky130_fd_sc_hd__dfxtp_2
X_11657_ _13721_/A1 hold1631/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11657_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12626__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13221__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12936__B1 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10608_ _10605_/Y _10788_/A _11596_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _10788_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14376_ _15441_/CLK _14376_/D vssd1 vssd1 vccd1 vccd1 _14376_/Q sky130_fd_sc_hd__dfxtp_1
X_11588_ _11588_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10947__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09000__A _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13327_ input149/X fanout5/X fanout3/X input117/X vssd1 vssd1 vccd1 vccd1 _13327_/X
+ sky130_fd_sc_hd__a22o_1
Xhold908 hold908/A vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ _10364_/X _10366_/Y _10537_/X _10538_/Y vssd1 vssd1 vccd1 vccd1 _10677_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold919 hold919/A vssd1 vssd1 vccd1 vccd1 hold919/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13258_ input156/X fanout6/X fanout4/X input124/X vssd1 vssd1 vccd1 vccd1 _13258_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08907__A2 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12209_ _14330_/Q _14234_/Q hold591/A hold985/A _12198_/S _12211_/S1 vssd1 vssd1
+ vccd1 vccd1 _12210_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _13393_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _15054_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2309 _06935_/Y vssd1 vssd1 vccd1 vccd1 _07457_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09580__A2 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13176__B _13176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1608 _13702_/X vssd1 vssd1 vccd1 vccd1 _15408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1619 _14348_/Q vssd1 vssd1 vccd1 vccd1 hold1619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07750_ _13655_/A1 hold2137/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07750_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09670__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ hold403/X _13654_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold404/A sky130_fd_sc_hd__mux2_1
XANTENNA__13192__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ _09420_/A _09420_/B _09420_/C vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09351_ _14440_/Q _09350_/C _09350_/A vssd1 vssd1 vccd1 vccd1 _09352_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08302_ _08312_/A _08702_/B _08228_/D _08225_/X vssd1 vssd1 vccd1 vccd1 _08314_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _09661_/A _09979_/C vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__and2_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11143__C _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08233_ _10873_/A _09437_/A vssd1 vssd1 vccd1 vccd1 _08234_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08164_ _08164_/A _08240_/A _08164_/C vssd1 vssd1 vccd1 vccd1 _08164_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07115_ _07115_/A _13502_/A vssd1 vssd1 vccd1 vccd1 _07115_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08095_ _08095_/A _08095_/B _08095_/C vssd1 vssd1 vccd1 vccd1 _08097_/A sky130_fd_sc_hd__and3_1
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07046_ _13651_/A1 hold2103/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07046_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12155__A1 _14984_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12271__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2810 _14282_/Q vssd1 vssd1 vccd1 vccd1 hold2810/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2821 _15051_/Q vssd1 vssd1 vccd1 vccd1 hold2821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2832 _15299_/Q vssd1 vssd1 vccd1 vccd1 hold443/A sky130_fd_sc_hd__dlygate4sd3_1
X_08997_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout764_A _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2843 _15302_/Q vssd1 vssd1 vccd1 vccd1 hold2843/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2854 _15321_/Q vssd1 vssd1 vccd1 vccd1 hold2854/X sky130_fd_sc_hd__dlygate4sd3_1
X_07948_ hold2755/X input26/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13175_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_199_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10469__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12863__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07879_ _07879_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__and2_4
XANTENNA__08908__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09618_ _11474_/A2 _09616_/X _09617_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _09618_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10890_ _10887_/X _10888_/Y _10704_/B _10707_/B vssd1 vssd1 vccd1 vccd1 _10890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09549_ _09549_/A _09549_/B _09549_/C vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__and3_2
XFILLER_0_109_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ hold965/A _13936_/Q _12560_/S vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_108_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11511_ _11509_/A _11500_/X _11510_/X _11511_/C1 vssd1 vssd1 vccd1 vccd1 _11512_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ hold851/A _14241_/Q _12491_/S vssd1 vssd1 vccd1 vccd1 _12491_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_136_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13041__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ _15418_/CLK hold836/X vssd1 vssd1 vccd1 vccd1 hold835/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _11441_/B _11441_/C _11441_/A vssd1 vssd1 vccd1 vccd1 _11443_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08047__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08135__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12394__A1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ _11586_/A _11614_/A _11564_/B _11614_/B vssd1 vssd1 vccd1 vccd1 _11374_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14161_ _15062_/CLK hold646/X vssd1 vssd1 vccd1 vccd1 hold645/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10324_ _10324_/A _10324_/B _10324_/C vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13112_ _13129_/A hold115/X vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__and2_1
XFILLER_0_131_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _14105_/CLK hold238/X vssd1 vssd1 vccd1 vccd1 _14092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13043_ _13098_/S1 _13040_/X _13042_/X vssd1 vssd1 vccd1 vccd1 _13043_/X sky130_fd_sc_hd__a21o_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10255_/A1 _10248_/Y _10250_/Y _10252_/Y _10254_/Y vssd1 vssd1 vccd1 vccd1
+ _10255_/X sky130_fd_sc_hd__o32a_1
XANTENNA__07275__A _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09562__A2 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ _10185_/A _11536_/B _10185_/C _10185_/D vssd1 vssd1 vccd1 vccd1 _10186_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_206_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14994_ _15250_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 _14994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13945_ _15377_/CLK _13945_/D vssd1 vssd1 vccd1 vccd1 _13945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13216__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ _14731_/CLK _13876_/D vssd1 vssd1 vccd1 vccd1 _13876_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07214__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10880__A1 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ _13102_/A _12827_/B _12827_/C vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__and3_1
XANTENNA__10880__B2 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _15408_/Q _14543_/Q hold911/A hold863/A _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12758_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__C1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ hold1009/X _13663_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12689_ hold757/X _14217_/Q hold605/A _14471_/Q _12591_/S _12689_/S1 vssd1 vssd1
+ vccd1 vccd1 _12689_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ _15299_/CLK _14428_/D vssd1 vssd1 vccd1 vccd1 _14428_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11188__A2 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14359_ _14909_/CLK hold630/X vssd1 vssd1 vccd1 vccd1 hold629/A sky130_fd_sc_hd__dfxtp_1
Xhold705 hold705/A vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12790__S _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold716 hold716/A vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold727 hold727/A vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 hold738/A vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 hold749/A vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__A1 hold2548/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13187__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09384__B _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10604__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2106 _07515_/X vssd1 vssd1 vccd1 vccd1 _14140_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A1 _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2117 _13918_/Q vssd1 vssd1 vccd1 vccd1 hold2117/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10243__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__B2 _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08851_ _08851_/A _09346_/B _08851_/C vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__or3_1
Xhold2128 _11940_/X vssd1 vssd1 vccd1 vccd1 _14760_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2139 _14372_/Q vssd1 vssd1 vccd1 vccd1 hold2139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1405 _15280_/Q vssd1 vssd1 vccd1 vccd1 hold1405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _07795_/X vssd1 vssd1 vccd1 vccd1 _14410_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ hold841/X _13740_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold842/A sky130_fd_sc_hd__mux2_1
XFILLER_0_209_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1427 _14110_/Q vssd1 vssd1 vccd1 vccd1 hold1427/X sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ _09009_/A _09866_/B _08783_/C _08783_/D vssd1 vssd1 vccd1 vccd1 _08782_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__13637__A1 _08107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1438 _11779_/X vssd1 vssd1 vccd1 vccd1 _14604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1449 _14313_/Q vssd1 vssd1 vccd1 vccd1 hold1449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13634__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__B1 _13468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ hold931/X _13739_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold932/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12030__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ hold1211/X _13736_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 _07664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07124__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _09542_/A _09979_/B _11407_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _09539_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07595_ _13734_/A1 hold1203/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07595_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12965__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _09330_/Y _09331_/X _09195_/Y _09197_/Y vssd1 vssd1 vccd1 vccd1 _09335_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09265_ _10110_/A _09726_/B _09264_/C _09264_/D vssd1 vssd1 vccd1 vccd1 _09266_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout512_A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12266__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _08297_/B _08214_/C _08214_/A vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__a21oi_1
X_09196_ _09196_/A _09196_/B vssd1 vssd1 vccd1 vccd1 _09198_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12376__A1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08147_/A _08147_/B _08147_/C vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__and3_1
XFILLER_0_161_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09241__A1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A2 _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08078_ _08077_/B _08077_/C _08077_/A vssd1 vssd1 vccd1 vccd1 _08080_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout881_A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07029_ hold1301/X _13519_/A0 _07044_/S vssd1 vssd1 vccd1 vccd1 _07029_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09294__B _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12679__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10040_ _09881_/A _09881_/C _09881_/B vssd1 vssd1 vccd1 vccd1 _10042_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09544__A2 _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2640 _08112_/Y vssd1 vssd1 vccd1 vccd1 hold2640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2651 _14447_/Q vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2662 _14818_/Q vssd1 vssd1 vccd1 vccd1 hold2662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2673 _12024_/X vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2684 _14436_/Q vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2695 _15190_/Q vssd1 vssd1 vccd1 vccd1 hold2695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1950 _11770_/X vssd1 vssd1 vccd1 vccd1 _14595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1961 _14761_/Q vssd1 vssd1 vccd1 vccd1 hold1961/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1972 _07196_/X vssd1 vssd1 vccd1 vccd1 _14003_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ hold287/X _13680_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__mux2_1
Xhold1983 _14535_/Q vssd1 vssd1 vccd1 vccd1 hold1983/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11103__A2 _11102_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ hold1133/X _13730_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 _13730_/X sky130_fd_sc_hd__mux2_1
Xhold1994 _11902_/X vssd1 vssd1 vccd1 vccd1 _14723_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ hold651/A _13954_/Q hold575/A _13922_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _10943_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07034__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ hold1013/X _13661_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 _13661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10873_ _10873_/A _15224_/Q vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__and2_1
XFILLER_0_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15400_ _15400_/CLK hold200/X vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__dfxtp_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ _12674_/S1 _12609_/X _12611_/X vssd1 vssd1 vccd1 vccd1 _12612_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12603__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ _14452_/Q _13636_/B vssd1 vssd1 vccd1 vccd1 _13592_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08654__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _15422_/CLK _15331_/D vssd1 vssd1 vccd1 vccd1 _15331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12668_/A1 _12540_/X _12542_/X vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__a21o_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15262_ _15364_/CLK _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/Q sky130_fd_sc_hd__dfxtp_1
X_12474_ _13868_/Q _13996_/Q _13836_/Q _13804_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12474_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13013__C1 hold2774/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_91_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ _15080_/CLK _14213_/D vssd1 vssd1 vccd1 vccd1 _14213_/Q sky130_fd_sc_hd__dfxtp_1
X_11425_ _11577_/A _11596_/A _14968_/Q _14969_/Q vssd1 vssd1 vccd1 vccd1 _11574_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15193_ _15196_/CLK _15193_/D vssd1 vssd1 vccd1 vccd1 _15193_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_111_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ _15364_/CLK _14144_/D vssd1 vssd1 vccd1 vccd1 _14144_/Q sky130_fd_sc_hd__dfxtp_1
X_11356_ _11356_/A _11518_/A _11356_/C vssd1 vssd1 vccd1 vccd1 _11518_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_46_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07794__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__B1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _10306_/A _11606_/A _10306_/C _10306_/D vssd1 vssd1 vccd1 vccd1 _10307_/X
+ sky130_fd_sc_hd__a22o_1
X_14075_ _14077_/CLK _14075_/D vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_11287_ _11283_/X _11286_/X _11287_/S vssd1 vssd1 vccd1 vccd1 _11287_/X sky130_fd_sc_hd__mux2_2
XANTENNA__10424__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07209__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ _13101_/A _13026_/B vssd1 vssd1 vccd1 vccd1 _13027_/C sky130_fd_sc_hd__or2_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10238_ hold279/A hold297/A hold311/A _13982_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10238_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_184_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11954__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10169_ _10169_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__or2_1
XFILLER_0_206_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09299__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14977_ _15250_/CLK hold116/X vssd1 vssd1 vccd1 vccd1 _14977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09299__B2 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10797__C _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13928_ _15398_/CLK hold976/X vssd1 vssd1 vccd1 vccd1 hold975/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_164_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12785__S _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13859_ _15458_/CLK hold946/X vssd1 vssd1 vccd1 vccd1 hold945/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_44_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13470__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ _07862_/B _14060_/Q _07404_/A _15344_/Q _07379_/X vssd1 vssd1 vccd1 vccd1
+ _07381_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__A1 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10605__B2 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_179_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12086__A _14983_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09050_ _09049_/B _09049_/C _09049_/A vssd1 vssd1 vccd1 vccd1 _09050_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_59_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12358__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ _07986_/Y _07991_/Y _08000_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08002_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08657__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold502 hold502/A vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold513 hold513/A vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 hold524/A vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold535 hold535/A vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__C _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 hold546/A vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold557 hold557/A vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 hold568/A vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _11499_/B1 _09945_/Y _09947_/Y _09949_/Y _09951_/Y vssd1 vssd1 vccd1 vccd1
+ _09952_/X sky130_fd_sc_hd__o32a_1
Xhold579 hold579/A vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _09021_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__and2_1
XANTENNA__07119__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _09883_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09886_/C sky130_fd_sc_hd__or2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07537__A1 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12530__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _11653_/X vssd1 vssd1 vccd1 vccd1 _14456_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ _08948_/A _08833_/B _08725_/A vssd1 vssd1 vccd1 vccd1 _08834_/X sky130_fd_sc_hd__o21ba_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _14381_/Q vssd1 vssd1 vccd1 vccd1 hold1213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1224 _11663_/X vssd1 vssd1 vccd1 vccd1 _14466_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1235 _14169_/Q vssd1 vssd1 vccd1 vccd1 hold1235/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1246 _11790_/X vssd1 vssd1 vccd1 vccd1 _14615_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1257 _14639_/Q vssd1 vssd1 vccd1 vccd1 hold1257/X sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ hold597/A _13939_/Q _15440_/Q _13907_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08766_/B sky130_fd_sc_hd__mux4_1
XANTENNA_fanout462_A _12056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 _11887_/X vssd1 vssd1 vccd1 vccd1 _14709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1279 _14393_/Q vssd1 vssd1 vccd1 vccd1 hold1279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ hold415/X _13689_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold416/A sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08696_ _09164_/A _09709_/B _08697_/A vssd1 vssd1 vccd1 vccd1 _08696_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ hold2203/X _13719_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 _07647_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout727_A _14960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12046__A0 _12112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07789__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ _12329_/A hold1183/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07578_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09317_ _09317_/A _09317_/B _09317_/C vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__or3_1
XFILLER_0_193_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10509__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _10142_/A _10142_/B _10126_/B vssd1 vssd1 vccd1 vccd1 _09248_/X sky130_fd_sc_hd__and3_1
XFILLER_0_146_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12349__A1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _09178_/B _09178_/C _09178_/A vssd1 vssd1 vccd1 vccd1 _09179_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__08648__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _11209_/B _11209_/C _11209_/A vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12190_ _14906_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12190_/X sky130_fd_sc_hd__or2_1
X_11141_ _11580_/A _14970_/Q vssd1 vssd1 vccd1 vccd1 _11578_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10244__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07029__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _10887_/X _10889_/Y _11070_/X _11071_/Y vssd1 vssd1 vccd1 vccd1 _11076_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput100 in1[12] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07528__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput111 in1[22] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_1
Xinput122 in1[3] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_1
X_10023_ _10024_/A _10024_/B _10024_/C vssd1 vssd1 vccd1 vccd1 _10023_/Y sky130_fd_sc_hd__nor3_1
X_14900_ _14987_/CLK _14900_/D vssd1 vssd1 vccd1 vccd1 _14900_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10758__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput133 in2[13] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__clkbuf_2
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput144 in2[23] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__clkbuf_2
Xinput155 in2[4] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09244__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2470 _12085_/X vssd1 vssd1 vccd1 vccd1 _14854_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _14876_/CLK _14831_/D vssd1 vssd1 vccd1 vccd1 _14831_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2481 _14847_/Q vssd1 vssd1 vccd1 vccd1 hold2481/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2492 _12121_/X vssd1 vssd1 vccd1 vccd1 _14872_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07272__B _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1780 _07176_/X vssd1 vssd1 vccd1 vccd1 _13984_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1791 _14265_/Q vssd1 vssd1 vccd1 vccd1 hold1791/X sky130_fd_sc_hd__dlygate4sd3_1
X_14762_ _15438_/CLK _14762_/D vssd1 vssd1 vccd1 vccd1 _14762_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ hold1377/X _13663_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11974_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ hold1765/X _13746_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13713_/X sky130_fd_sc_hd__mux2_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _14451_/Q _11113_/C vssd1 vssd1 vccd1 vccd1 _10925_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_168_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14693_ _15398_/CLK hold816/X vssd1 vssd1 vccd1 vccd1 hold815/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11225__D _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13290__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07699__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13644_ input54/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13644_/X sky130_fd_sc_hd__or2_1
X_10856_ _11037_/A _10856_/B _10856_/C _10856_/D vssd1 vssd1 vccd1 vccd1 _11037_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12588__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _09625_/A _13586_/B _13574_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13575_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ _10787_/A _10787_/B vssd1 vssd1 vccd1 vccd1 _10790_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12683__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15315_/CLK _15314_/D vssd1 vssd1 vccd1 vccd1 _15314_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12526_ _12601_/A _12526_/B vssd1 vssd1 vccd1 vccd1 _12527_/C sky130_fd_sc_hd__or2_1
XFILLER_0_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11949__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _15247_/CLK hold122/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12457_ _12607_/A _12457_/B vssd1 vssd1 vccd1 vccd1 _14946_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11408_ _11408_/A _11408_/B vssd1 vssd1 vccd1 vccd1 _11410_/A sky130_fd_sc_hd__nor2_1
X_15176_ _15177_/CLK _15176_/D vssd1 vssd1 vccd1 vccd1 _15176_/Q sky130_fd_sc_hd__dfxtp_1
X_12388_ _12642_/B1 _12383_/X _12387_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12395_/A
+ sky130_fd_sc_hd__o211a_1
X_14127_ _15448_/CLK _14127_/D vssd1 vssd1 vccd1 vccd1 _14127_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07447__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11339_ _11339_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10154__A _10154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09943__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14058_ _15351_/CLK _14058_/D vssd1 vssd1 vccd1 vccd1 hold573/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12512__A1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11684__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09913__C1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ hold575/X hold2135/X _13041_/S vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13184__B _13184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08550_ _08197_/A _08547_/X _08549_/X vssd1 vssd1 vccd1 vccd1 _08550_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09367__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07501_ hold2043/X _13740_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07501_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12371__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08481_ _08480_/B _08480_/C _08480_/A vssd1 vssd1 vccd1 vccd1 _08483_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12028__A0 hold2562/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07432_ _07432_/A _07450_/B vssd1 vssd1 vccd1 vccd1 _14062_/D sky130_fd_sc_hd__and2_1
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08294__A _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07363_ _13081_/A1 _07904_/B _14022_/Q vssd1 vssd1 vccd1 vccd1 _12308_/A sky130_fd_sc_hd__a21boi_2
XANTENNA_hold2859_A _15341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12674__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ _09514_/A _09099_/X _09101_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09103_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07294_ _15223_/Q _14967_/Q vssd1 vssd1 vccd1 vccd1 _07296_/A sky130_fd_sc_hd__or2_1
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13528__A0 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11859__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12263__B _13412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold332 hold332/A vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 hold343/A vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold365 hold365/A vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 hold376/A vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold387 hold387/A vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 hold398/A vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _12689_/S1 vssd1 vssd1 vccd1 vccd1 _12474_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout812 _12939_/S1 vssd1 vssd1 vccd1 vccd1 _12949_/S1 sky130_fd_sc_hd__clkbuf_8
X_09935_ hold205/A hold559/A hold507/A _13980_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _09935_/X sky130_fd_sc_hd__mux4_1
Xfanout823 _12641_/S vssd1 vssd1 vccd1 vccd1 _12441_/S sky130_fd_sc_hd__buf_8
Xfanout834 _12915_/S vssd1 vssd1 vccd1 vccd1 _12916_/S sky130_fd_sc_hd__buf_8
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13375__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _13178_/A vssd1 vssd1 vccd1 vccd1 _13565_/C1 sky130_fd_sc_hd__buf_4
Xfanout856 _13535_/B vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__clkbuf_4
X_09866_ _10022_/B _09866_/B _09866_/C _09866_/D vssd1 vssd1 vccd1 vccd1 _09869_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 _13490_/A vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__buf_2
Xfanout878 _13479_/A vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08469__A _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 _11709_/X vssd1 vssd1 vccd1 vccd1 _14505_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1021 _15075_/Q vssd1 vssd1 vccd1 vccd1 hold1021/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 _13338_/A vssd1 vssd1 vccd1 vccd1 _13390_/A sky130_fd_sc_hd__buf_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _08820_/B vssd1 vssd1 vccd1 vccd1 _08817_/Y sky130_fd_sc_hd__inv_2
Xhold1032 _13215_/X vssd1 vssd1 vccd1 vccd1 _15079_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _15263_/Q vssd1 vssd1 vccd1 vccd1 hold1043/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout844_A _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ hold979/A _14223_/Q hold389/A _14477_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09798_/B sky130_fd_sc_hd__mux4_1
Xhold1054 _11968_/X vssd1 vssd1 vccd1 vccd1 _14787_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07930__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 _14151_/Q vssd1 vssd1 vccd1 vccd1 hold1065/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 _13481_/X vssd1 vssd1 vccd1 vccd1 _15240_/D sky130_fd_sc_hd__buf_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09358__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _09918_/A _13430_/B _08747_/X _10233_/A vssd1 vssd1 vccd1 vccd1 _08748_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1087 _14746_/Q vssd1 vssd1 vccd1 vccd1 hold1087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12806__A2 _13159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_205 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1098 _13209_/X vssd1 vssd1 vccd1 vccd1 _15073_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_216 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12362__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08678_/B _08678_/C _08678_/A vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10710_ _10706_/X _10708_/Y _10532_/B _10534_/B vssd1 vssd1 vccd1 vccd1 _10710_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11623__A _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _06905_/A _13792_/A2 _11689_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _14490_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__and2_1
XFILLER_0_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13360_ _13360_/A _13360_/B vssd1 vssd1 vccd1 vccd1 _15151_/D sky130_fd_sc_hd__nor2_1
X_10572_ _13586_/A _10571_/B _10751_/B _10233_/A vssd1 vssd1 vccd1 vccd1 _10572_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_180_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11769__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ _14330_/Q _14234_/Q hold591/A hold985/A _12365_/S0 _12365_/S1 vssd1 vssd1
+ vccd1 vccd1 _12311_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13291_ input136/X fanout5/X fanout3/X input104/X vssd1 vssd1 vccd1 vccd1 _13291_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _15190_/CLK _15030_/D vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07548__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _14331_/Q _14235_/Q _14395_/Q hold895/A _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12243_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12742__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ hold2591/X _12173_/A2 _12172_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ hold287/A hold413/A hold727/A _14746_/Q _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _11125_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_120_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11055_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__xor2_1
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10006_ _10115_/A _10283_/C _10115_/D _10110_/A vssd1 vssd1 vccd1 vccd1 _10010_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11517__B _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14814_ _14844_/CLK _14814_/D vssd1 vssd1 vccd1 vccd1 _14814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09123__B1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _15421_/CLK _14745_/D vssd1 vssd1 vccd1 vccd1 _14745_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ hold2809/X hold1629/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11957_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09674__A1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09674__B2 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13224__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ _10690_/X _10693_/Y _11098_/A _10907_/X vssd1 vssd1 vccd1 vccd1 _11098_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__10284__A2 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14676_ _15450_/CLK hold608/X vssd1 vssd1 vccd1 vccd1 hold607/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11888_ hold331/X _13742_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold332/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ hold2569/X _13797_/A2 _13626_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15341_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08229__A2 _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ _11570_/A _11537_/A _11623_/B _11605_/A vssd1 vssd1 vccd1 vccd1 _10840_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09977__A2 _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ _13558_/A _13570_/B vssd1 vssd1 vccd1 vccd1 _13558_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12981__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ _15435_/Q _13902_/Q _12566_/S vssd1 vssd1 vccd1 vccd1 _12509_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09657__B _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ _13489_/A hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__and2_1
XFILLER_0_180_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12408__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15228_ _15324_/CLK _15228_/D vssd1 vssd1 vccd1 vccd1 _15228_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10419__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15159_ _15320_/CLK _15159_/D vssd1 vssd1 vccd1 vccd1 _15159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07981_ _07981_/A _07981_/B _07981_/C vssd1 vssd1 vccd1 vccd1 _07981_/X sky130_fd_sc_hd__or3_1
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09720_ _09720_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__13195__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06932_ _14088_/Q vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__inv_2
XFILLER_0_207_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11427__B _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _09636_/Y _09641_/Y _09650_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09652_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08602_ _09138_/A _08809_/B _08809_/D _08776_/B vssd1 vssd1 vccd1 vccd1 _08604_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12249__B1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09582_ _10110_/A _10115_/A _09724_/C _09724_/D vssd1 vssd1 vccd1 vccd1 _09584_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_171_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08533_ _07900_/B _08532_/Y _08467_/X vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13461__A2 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10985__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08464_ _08449_/Y _08454_/Y _08463_/X _12241_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08465_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07132__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07415_ hold95/X _07448_/B vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__and2_1
XFILLER_0_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08395_ _09816_/A _08685_/C _08395_/C _08395_/D vssd1 vssd1 vccd1 vccd1 _08397_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12647__S1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_A _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11224__A1 _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__B2 _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ _07346_/A _15332_/Q vssd1 vssd1 vccd1 vccd1 _07362_/C sky130_fd_sc_hd__or2_1
XFILLER_0_190_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10432__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07277_ _09075_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07327_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12274__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09016_ _09016_/A _09016_/B vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13072__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout620 _10142_/A vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__clkbuf_8
Xfanout631 _15202_/Q vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__clkbuf_4
Xfanout642 _08075_/B vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__buf_2
X_09918_ _09918_/A _13448_/B vssd1 vssd1 vccd1 vccd1 _09918_/Y sky130_fd_sc_hd__nor2_1
Xfanout653 _15197_/Q vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08199__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 _15063_/Q vssd1 vssd1 vccd1 vccd1 _13743_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout675 _13705_/A1 vssd1 vssd1 vccd1 vccd1 _13738_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__09353__B1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout686 _13700_/A1 vssd1 vssd1 vccd1 vccd1 _13519_/A0 sky130_fd_sc_hd__clkbuf_4
X_09849_ _10110_/A _10283_/C _10115_/D _10002_/C vssd1 vssd1 vccd1 vccd1 _09851_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10879__D _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout697 _15048_/Q vssd1 vssd1 vccd1 vccd1 _13662_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_198_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ hold445/A _13948_/Q _13066_/S vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__mux2_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12335__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ hold887/X _13665_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold888/A sky130_fd_sc_hd__mux2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _14349_/Q _14253_/Q _12791_/S vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__mux2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14530_ _15432_/CLK _14530_/D vssd1 vssd1 vccd1 vccd1 _14530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _13728_/A1 hold2177/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11742_/X sky130_fd_sc_hd__mux2_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07042__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ _14754_/CLK _14461_/D vssd1 vssd1 vccd1 vccd1 _14461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11673_ _13704_/A1 hold1763/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10018__A2 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ _13450_/A _13412_/B vssd1 vssd1 vccd1 vccd1 _13412_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09959__A2 _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10624_ _11590_/A _11605_/B _10623_/C _10623_/D vssd1 vssd1 vccd1 vccd1 _10624_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ _15457_/CLK _14392_/D vssd1 vssd1 vccd1 vccd1 _14392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08662__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12963__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11310__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ _13369_/A _13343_/B vssd1 vssd1 vccd1 vccd1 _15134_/D sky130_fd_sc_hd__nor2_1
X_10555_ _10382_/Y _10387_/A _10553_/X _10554_/Y vssd1 vssd1 vccd1 vccd1 _10557_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07278__A _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ input66/X fanout1/X _13273_/X vssd1 vssd1 vccd1 vccd1 _13275_/B sky130_fd_sc_hd__a21oi_1
X_10486_ _11569_/A _11537_/A _11623_/B _11563_/A vssd1 vssd1 vccd1 vccd1 _10487_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output177_A _15188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15013_ _15179_/CLK _15013_/D vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12225_ _07900_/B _12223_/Y _13172_/B _12259_/A1 _12219_/X vssd1 vssd1 vccd1 vccd1
+ _12225_/X sky130_fd_sc_hd__a221o_1
X_12156_ _12156_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13219__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _11107_/A _11481_/A vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__nand2_1
X_12087_ hold2457/X _12129_/A2 _12086_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12087_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12574__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ _10893_/B _11038_/B vssd1 vssd1 vccd1 vccd1 _11081_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__11247__B _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12745__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ hold1861/X hold1597/X hold633/X hold1513/X _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12989_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_176_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14728_ _15268_/CLK _14728_/D vssd1 vssd1 vccd1 vccd1 _14728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12895__C_N _13076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14659_ _14754_/CLK hold466/X vssd1 vssd1 vccd1 vccd1 _14659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_180_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15434_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07200_ hold291/X _13668_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__mux2_1
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10009__A2 _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12403__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ _08178_/Y _08180_/B vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08572__A _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12954__A1 _10566_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ _13732_/A1 hold2019/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07131_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11301__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2557_A _15352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__A _14987_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08291__B _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07062_ _13519_/A0 hold1789/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07062_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput201 _14184_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[14] sky130_fd_sc_hd__buf_12
XFILLER_0_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12706__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput212 _14194_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[24] sky130_fd_sc_hd__buf_12
XFILLER_0_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput223 _14175_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[5] sky130_fd_sc_hd__buf_12
Xoutput234 _14439_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[15] sky130_fd_sc_hd__buf_12
XFILLER_0_65_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput245 _14449_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[25] sky130_fd_sc_hd__buf_12
Xoutput256 _14430_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[6] sky130_fd_sc_hd__buf_12
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4__f_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput267 _14893_/Q vssd1 vssd1 vccd1 vccd1 out0[16] sky130_fd_sc_hd__buf_12
XFILLER_0_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput278 _14903_/Q vssd1 vssd1 vccd1 vccd1 out0[26] sky130_fd_sc_hd__buf_12
XFILLER_0_11_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput289 _14884_/Q vssd1 vssd1 vccd1 vccd1 out0[7] sky130_fd_sc_hd__buf_12
XFILLER_0_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11438__A _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07964_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07964_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09703_ _10110_/A _10010_/B _09700_/Y _09701_/X vssd1 vssd1 vccd1 vccd1 _09704_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07127__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ _14446_/Q vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__inv_2
XFILLER_0_208_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07895_ _07895_/A vssd1 vssd1 vccd1 vccd1 _07965_/A sky130_fd_sc_hd__inv_2
XANTENNA__11142__B1 _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11872__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _13502_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _13882_/Q hold617/A hold659/A _13818_/Q _10425_/S0 _10425_/S1 vssd1 vssd1
+ vccd1 vccd1 _09634_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09850__B _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__B1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13419__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12317__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09565_ _10129_/A _11407_/A vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout542_A _15423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _08516_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12642__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ _13590_/B _09494_/Y _09495_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _09496_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ _13872_/Q _14000_/Q _13840_/Q _13808_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08447_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_171_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15371_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout807_A _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ _08378_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08378_/X sky130_fd_sc_hd__or2_1
XFILLER_0_191_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07329_ _12254_/B _07329_/B _07329_/C _07328_/X vssd1 vssd1 vccd1 vccd1 _07330_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_116_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__B _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10340_ _10338_/X _10340_/B vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _11580_/A _11578_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _10273_/B sky130_fd_sc_hd__and3_1
XFILLER_0_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ hold2621/X hold2662/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07826__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__A1 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10184__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10252__A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 _07981_/A vssd1 vssd1 vccd1 vccd1 _13554_/B sky130_fd_sc_hd__clkbuf_2
Xfanout461 _12062_/S vssd1 vssd1 vccd1 vccd1 _12058_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__07037__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout472 _08637_/Y vssd1 vssd1 vccd1 vccd1 _13031_/B1 sky130_fd_sc_hd__buf_4
X_13961_ _15072_/CLK _13961_/D vssd1 vssd1 vccd1 vccd1 _13961_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09877__A1 _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout483 _07862_/X vssd1 vssd1 vccd1 vccd1 _11511_/C1 sky130_fd_sc_hd__buf_8
Xfanout494 _06944_/Y vssd1 vssd1 vccd1 vccd1 _13100_/S1 sky130_fd_sc_hd__buf_8
XANTENNA__11782__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _12949_/S1 _12909_/X _12911_/X vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _14651_/CLK _13892_/D vssd1 vssd1 vccd1 vccd1 _13892_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12881__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ _12939_/S1 _12840_/X _12842_/X vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__a21o_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_15__f_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ _13880_/Q _14008_/Q hold663/A _13816_/Q _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12774_/X sky130_fd_sc_hd__mux4_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _15376_/CLK _14513_/D vssd1 vssd1 vccd1 vccd1 _14513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ hold349/X _13679_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 hold350/A sky130_fd_sc_hd__mux2_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_162_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14444_ _15316_/CLK _14444_/D vssd1 vssd1 vccd1 vccd1 _14444_/Q sky130_fd_sc_hd__dfxtp_1
X_11656_ _13687_/A1 hold1981/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11656_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07500__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12936__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _11596_/A _11594_/B _10605_/Y _10788_/A vssd1 vssd1 vccd1 vccd1 _10609_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14375_ _15371_/CLK _14375_/D vssd1 vssd1 vccd1 vccd1 _14375_/Q sky130_fd_sc_hd__dfxtp_1
X_11587_ _11587_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ _13338_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _15128_/D sky130_fd_sc_hd__nor2_1
X_10538_ _10534_/X _10535_/Y _10362_/B _10364_/B vssd1 vssd1 vccd1 vccd1 _10538_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10411__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold909 hold909/A vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11957__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ _13287_/A _13257_/B vssd1 vssd1 vccd1 vccd1 _15105_/D sky130_fd_sc_hd__nor2_1
X_10469_ _11614_/A _10827_/D _11537_/B _11586_/A vssd1 vssd1 vccd1 vccd1 _10469_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _12241_/A _12208_/B _12208_/C vssd1 vssd1 vccd1 vccd1 _12219_/C sky130_fd_sc_hd__or3_1
XFILLER_0_209_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13188_ _13396_/A _13188_/B vssd1 vssd1 vccd1 vccd1 _15053_/D sky130_fd_sc_hd__and2_1
XFILLER_0_202_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11372__B1 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ hold2586/X _12195_/A2 _12138_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12139_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13649__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1609 _15288_/Q vssd1 vssd1 vccd1 vccd1 hold1609/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12547__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13473__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__B _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__A2 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ hold301/X _13653_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__mux2_1
XANTENNA__08540__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09350_ _09350_/A _09350_/B _09350_/C vssd1 vssd1 vccd1 vccd1 _09498_/C sky130_fd_sc_hd__and3_1
XFILLER_0_133_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08301_ _08301_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _09816_/A _09979_/D vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__nand2_1
XANTENNA_hold2674_A _14828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11143__D _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_153_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15367_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08234_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12388__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _08162_/A _08162_/B _08162_/C vssd1 vssd1 vccd1 vccd1 _08164_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12028__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07114_ _14087_/Q _07114_/B vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__or2_4
X_08094_ _08093_/A _08093_/B _08093_/C vssd1 vssd1 vccd1 vccd1 _08095_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11867__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13648__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07045_ _14086_/Q _14087_/Q _07182_/A _07643_/C vssd1 vssd1 vccd1 vccd1 _07045_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout492_A _06944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2800 _15414_/Q vssd1 vssd1 vccd1 vccd1 hold2800/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2811 _14706_/Q vssd1 vssd1 vccd1 vccd1 hold2811/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08996_ _13732_/A1 _11514_/A2 _11514_/B1 _13187_/B _08994_/Y vssd1 vssd1 vccd1 vccd1
+ _08996_/X sky130_fd_sc_hd__a221o_1
Xhold2822 _15049_/Q vssd1 vssd1 vccd1 vccd1 hold2822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2833 _15306_/Q vssd1 vssd1 vccd1 vccd1 hold2833/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13104__A1 _11641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2844 _15298_/Q vssd1 vssd1 vccd1 vccd1 hold2844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2855 _14455_/Q vssd1 vssd1 vccd1 vccd1 hold2855/X sky130_fd_sc_hd__dlygate4sd3_1
X_07947_ _12252_/B _07947_/B vssd1 vssd1 vccd1 vccd1 _07947_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_199_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09859__A1 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10469__A2 _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _12301_/A _07878_/B _07878_/C _07846_/A vssd1 vssd1 vccd1 vccd1 _07899_/A
+ sky130_fd_sc_hd__or4b_4
XANTENNA__08477__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08908__C _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _09617_/A _11283_/S vssd1 vssd1 vccd1 vccd1 _09617_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13407__A2 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ _09547_/B _09547_/C _09547_/A vssd1 vssd1 vccd1 vccd1 _09549_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12431__A1_N _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09479_ _09478_/A _09478_/B _10397_/A vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_148_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_144_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15287_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12727__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _11510_/A1 _11502_/Y _11504_/Y _11509_/Y vssd1 vssd1 vccd1 vccd1 _11510_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12490_ hold441/X _14113_/Q _12491_/S vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09101__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12918__A1 _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _11441_/A _11441_/B _11441_/C vssd1 vssd1 vccd1 vccd1 _11443_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_163_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14160_ _15380_/CLK hold692/X vssd1 vssd1 vccd1 vccd1 hold691/A sky130_fd_sc_hd__dfxtp_1
X_11372_ _11614_/A _11564_/B _11614_/B _11586_/A vssd1 vssd1 vccd1 vccd1 _11374_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11777__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ _13129_/A hold61/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__and2_1
X_10323_ _10324_/A _10324_/B _10324_/C vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__and3_1
X_14091_ _14105_/CLK _14091_/D vssd1 vssd1 vccd1 vccd1 _14091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _13092_/A1 _13041_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07556__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ _15424_/Q _10253_/X _10255_/A1 vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09642__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10185_ _10185_/A _11378_/D _10185_/C _10185_/D vssd1 vssd1 vccd1 vccd1 _10185_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08770__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14993_ _15250_/CLK hold138/X vssd1 vssd1 vccd1 vccd1 _14993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13293__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13944_ _15408_/CLK _13944_/D vssd1 vssd1 vccd1 vccd1 _13944_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08387__A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07291__A _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ _15369_/CLK _13875_/D vssd1 vssd1 vccd1 vccd1 _13875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12826_ _12951_/A _12826_/B vssd1 vssd1 vccd1 vccd1 _12827_/C sky130_fd_sc_hd__or2_1
XANTENNA__10880__A2 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12606__B1 _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12757_ _13107_/A _12757_/B vssd1 vssd1 vccd1 vccd1 _14958_/D sky130_fd_sc_hd__nor2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_135_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15450_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11541__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11708_ hold1651/X _13662_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11708_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ _12366_/A _12683_/X _12687_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12695_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14427_ _15304_/CLK _14427_/D vssd1 vssd1 vccd1 vccd1 _14427_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11639_ _11469_/Y _11473_/C _11637_/Y _11638_/Y _08526_/B vssd1 vssd1 vccd1 vccd1
+ _11639_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13031__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14358_ _14485_/CLK _14358_/D vssd1 vssd1 vccd1 vccd1 _14358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 hold706/A vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 hold717/A vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ input143/X fanout5/X fanout3/X input111/X vssd1 vssd1 vccd1 vccd1 _13309_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13468__A _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 hold728/A vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold739 hold739/A vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ _15450_/CLK _14289_/D vssd1 vssd1 vccd1 vccd1 _14289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09633__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__B _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2107 _14513_/Q vssd1 vssd1 vccd1 vccd1 hold2107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _09346_/B _08851_/C _08851_/A vssd1 vssd1 vccd1 vccd1 _08850_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10699__A2 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2118 _07105_/X vssd1 vssd1 vccd1 vccd1 _13918_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10243__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2129 _14740_/Q vssd1 vssd1 vccd1 vccd1 hold2129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1406 _13522_/X vssd1 vssd1 vccd1 vccd1 _15280_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07801_ hold501/X _13739_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold502/A sky130_fd_sc_hd__mux2_1
X_08781_ _08901_/A _08892_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _08783_/D
+ sky130_fd_sc_hd__nand4_1
Xhold1417 _15269_/Q vssd1 vssd1 vccd1 vccd1 hold1417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 _07482_/X vssd1 vssd1 vccd1 vccd1 _14110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1439 _14770_/Q vssd1 vssd1 vccd1 vccd1 hold1439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11648__A1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ hold383/X _13738_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold384/A sky130_fd_sc_hd__mux2_1
XANTENNA__11648__B2 _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07663_ hold673/X _15055_/Q _07676_/S vssd1 vssd1 vccd1 vccd1 hold674/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09402_ _09979_/B _11407_/A _15209_/Q _10183_/A vssd1 vssd1 vccd1 vccd1 _09404_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07594_ _13700_/A1 hold1011/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07594_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09333_ _09330_/Y _09331_/X _09195_/Y _09197_/Y vssd1 vssd1 vccd1 vccd1 _09333_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_126_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15444_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10084__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ _10110_/A _09726_/B _09264_/C _09264_/D vssd1 vssd1 vccd1 vccd1 _09449_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07140__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _08301_/A vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__inv_2
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09195_ _09196_/A _09196_/B vssd1 vssd1 vccd1 vccd1 _09195_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout505_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08124__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _08077_/A _08077_/C _08077_/B vssd1 vssd1 vccd1 vccd1 _08147_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08760__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13378__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ _08077_/A _08077_/B _08077_/C vssd1 vssd1 vccd1 vccd1 _08080_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12282__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13325__A1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07028_ hold1769/X _13666_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout874_A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11887__A1 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2630 _14443_/Q vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2641 _15344_/Q vssd1 vssd1 vccd1 vccd1 hold2641/X sky130_fd_sc_hd__buf_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ hold845/A hold947/A _15084_/Q _14377_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _08979_/X sky130_fd_sc_hd__mux4_1
Xhold2652 _10237_/X vssd1 vssd1 vccd1 vccd1 _14447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2663 _14440_/Q vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08919__B _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2674 _14828_/Q vssd1 vssd1 vccd1 vccd1 hold2674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1940 _11969_/X vssd1 vssd1 vccd1 vccd1 _14788_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2685 _08751_/X vssd1 vssd1 vccd1 vccd1 _14436_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1951 _14736_/Q vssd1 vssd1 vccd1 vccd1 hold1951/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2696 _14844_/Q vssd1 vssd1 vccd1 vccd1 hold2696/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12836__B1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11990_ hold371/X _13679_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__mux2_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1962 _11941_/X vssd1 vssd1 vccd1 vccd1 _14761_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1973 _14065_/Q vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1984 _11741_/X vssd1 vssd1 vccd1 vccd1 _14535_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11345__B _15227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1995 _14297_/Q vssd1 vssd1 vccd1 vccd1 hold1995/X sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _11504_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ hold339/X _13693_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold340/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _10872_/A _10872_/B vssd1 vssd1 vccd1 vccd1 _10875_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12642_/A1 _12610_/X _12700_/S0 vssd1 vssd1 vccd1 vccd1 _12611_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13560__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08268__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_117_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15087_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11498__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ _10921_/B _13591_/A2 _13590_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _15321_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15340_/CLK _15330_/D vssd1 vssd1 vccd1 vccd1 _15330_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12692_/A1 _12541_/X _14490_/Q vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07050__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15261_ _15261_/CLK _15261_/D vssd1 vssd1 vccd1 vccd1 _15261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12473_ hold187/A hold333/A _14595_/Q _13964_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12473_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12891__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14212_ _15437_/CLK _14212_/D vssd1 vssd1 vccd1 vccd1 _14212_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08115__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11424_ _11596_/A _14968_/Q _14969_/Q _11577_/A vssd1 vssd1 vccd1 vccd1 _11427_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _15196_/CLK _15192_/D vssd1 vssd1 vccd1 vccd1 _15192_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__08670__A _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14143_ _14754_/CLK _14143_/D vssd1 vssd1 vccd1 vccd1 _14143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _11354_/B _11354_/C _11354_/A vssd1 vssd1 vccd1 vccd1 _11356_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__A1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ _10306_/A _11606_/A _10306_/C _10306_/D vssd1 vssd1 vccd1 vccd1 _10306_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__07286__A _15228_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14074_ _14077_/CLK _14074_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
X_11286_ _11286_/A _11286_/B vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output257_A _14431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ _13021_/X _13022_/X _13024_/X _13023_/X _13050_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _13026_/B sky130_fd_sc_hd__mux4_1
X_10237_ _10232_/A _13797_/A2 _10236_/Y _13797_/C1 vssd1 vssd1 vccd1 vccd1 _10237_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10168_ _10165_/Y _10343_/A _11335_/A _10338_/D vssd1 vssd1 vccd1 vccd1 _10343_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11536__A _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13227__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09299__A2 _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14976_ _15250_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 _14976_/Q sky130_fd_sc_hd__dfxtp_1
X_10099_ hold607/A _13949_/Q hold329/A _13917_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10100_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_178_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07929__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__D _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ _15428_/CLK _13927_/D vssd1 vssd1 vccd1 vccd1 _13927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10302__A1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10302__B2 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11970__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13858_ _15196_/CLK _13858_/D vssd1 vssd1 vccd1 vccd1 _13858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12809_ hold915/X _13914_/Q _12841_/S vssd1 vssd1 vccd1 vccd1 _12809_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15378_/CLK sky130_fd_sc_hd__clkbuf_16
X_13789_ _13241_/A _13625_/C _11687_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _15347_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10605__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12086__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15459_ _15460_/CLK _15459_/D vssd1 vssd1 vccd1 vccd1 _15459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08000_ _08564_/A1 _07993_/Y _07995_/Y _07997_/Y _07999_/Y vssd1 vssd1 vccd1 vccd1
+ _08000_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_154_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09676__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12989__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08657__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12763__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 hold503/A vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13198__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 hold525/A vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold536 hold536/A vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__D _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold547 hold547/A vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08982__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 hold558/A vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _11507_/A _09950_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _09951_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold569 hold569/A vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ _08901_/A _09726_/B _08901_/C vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _09881_/B _09881_/C _09881_/A vssd1 vssd1 vccd1 vccd1 _09883_/B sky130_fd_sc_hd__a21oi_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ _08948_/A _08833_/B _08725_/A vssd1 vssd1 vccd1 vccd1 _08953_/A sky130_fd_sc_hd__nor3b_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _14219_/Q vssd1 vssd1 vccd1 vccd1 hold1203/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _07765_/X vssd1 vssd1 vccd1 vccd1 _14381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 _14515_/Q vssd1 vssd1 vccd1 vccd1 hold1225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1236 _07544_/X vssd1 vssd1 vccd1 vccd1 _14169_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08989_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08764_/Y sky130_fd_sc_hd__nor2_1
Xhold1247 _14668_/Q vssd1 vssd1 vccd1 vccd1 hold1247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 _11815_/X vssd1 vssd1 vccd1 vccd1 _14639_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1269 _15436_/Q vssd1 vssd1 vccd1 vccd1 hold1269/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ hold603/X _13721_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold604/A sky130_fd_sc_hd__mux2_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _09164_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _08697_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout455_A _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11880__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ hold509/X _13718_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold510/A sky130_fd_sc_hd__mux2_1
XFILLER_0_138_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13380__B _13380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07577_ _13502_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _07577_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_165_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout622_A _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12277__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09316_ _09317_/A _09317_/B _09317_/C vssd1 vssd1 vccd1 vccd1 _09316_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_192_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__B _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09247_ _10142_/B _10126_/A _10126_/B _10142_/A vssd1 vssd1 vccd1 vccd1 _09247_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09178_ _09178_/A _09178_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09178_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08648__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ _08201_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11140_ _13746_/A1 _11514_/A2 _11514_/B1 _13201_/B _11138_/Y vssd1 vssd1 vccd1 vccd1
+ _11140_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11071_ _11067_/X _11068_/Y _10885_/B _10887_/B vssd1 vssd1 vccd1 vccd1 _11071_/Y
+ sky130_fd_sc_hd__o211ai_2
Xinput101 in1[13] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08186__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput112 in1[23] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10022_ _10022_/A _10022_/B _10304_/C _10304_/D vssd1 vssd1 vccd1 vccd1 _10024_/C
+ sky130_fd_sc_hd__and4_1
Xinput123 in1[4] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_1
Xinput134 in2[14] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__clkbuf_2
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 in2[24] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__clkbuf_2
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2460 _12115_/X vssd1 vssd1 vccd1 vccd1 _14869_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput156 in2[5] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _14866_/CLK _14830_/D vssd1 vssd1 vccd1 vccd1 _14830_/Q sky130_fd_sc_hd__dfxtp_2
Xhold2471 _14989_/Q vssd1 vssd1 vccd1 vccd1 hold2471/X sky130_fd_sc_hd__clkbuf_2
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2482 _12071_/X vssd1 vssd1 vccd1 vccd1 _14847_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2493 _14871_/Q vssd1 vssd1 vccd1 vccd1 hold2493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1770 _07028_/X vssd1 vssd1 vccd1 vccd1 _13845_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11973_ hold1605/X _13662_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__mux2_1
X_14761_ _15440_/CLK _14761_/D vssd1 vssd1 vccd1 vccd1 _14761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1781 _14388_/Q vssd1 vssd1 vccd1 vccd1 hold1781/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1792 _07642_/X vssd1 vssd1 vccd1 vccd1 _14265_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11790__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ hold807/X _13745_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold808/A sky130_fd_sc_hd__mux2_1
X_10924_ _13750_/A _13369_/B vssd1 vssd1 vccd1 vccd1 _10924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_169_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _15397_/CLK hold544/X vssd1 vssd1 vccd1 vccd1 hold543/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _08345_/A _13625_/C _13642_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15354_/D
+ sky130_fd_sc_hd__o211a_1
X_10855_ _10852_/X _10853_/Y _10663_/X _10668_/A vssd1 vssd1 vccd1 vccd1 _10856_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _14443_/Q _13590_/B vssd1 vssd1 vccd1 vccd1 _13574_/X sky130_fd_sc_hd__or2_1
X_10786_ _11597_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _10787_/B sky130_fd_sc_hd__nand2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _15313_/CLK _15313_/D vssd1 vssd1 vccd1 vccd1 _15313_/Q sky130_fd_sc_hd__dfxtp_1
X_12525_ _12521_/X _12522_/X _12524_/X _12523_/X _12669_/A1 _12700_/S1 vssd1 vssd1
+ vccd1 vccd1 _12526_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13510__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12456_ _08107_/A _08636_/A _13145_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12457_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ _15244_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11407_ _11407_/A _11570_/A _11606_/B _11570_/B vssd1 vssd1 vccd1 vccd1 _11408_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15175_ _15177_/CLK _15175_/D vssd1 vssd1 vccd1 vccd1 _15175_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ _12599_/S1 _12384_/X _12386_/X vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14126_ _15089_/CLK hold942/X vssd1 vssd1 vccd1 vccd1 hold941/A sky130_fd_sc_hd__dfxtp_1
X_11338_ _11339_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11338_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11965__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _15351_/CLK _14057_/D vssd1 vssd1 vccd1 vccd1 _14057_/Q sky130_fd_sc_hd__dfxtp_1
X_11269_ _11465_/A _11269_/B _11269_/C vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ hold807/X hold1491/X hold731/X hold1629/X _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13008_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_20_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14959_ _14971_/CLK _14959_/D vssd1 vssd1 vccd1 vccd1 _14959_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13481__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ hold1671/X _13739_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07500_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_159_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08480_ _08480_/A _08480_/B _08480_/C vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12371__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07431_ _07431_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14061_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08294__B _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12579__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07362_ _07427_/A _07362_/B _07362_/C _07362_/D vssd1 vssd1 vccd1 vccd1 _07904_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_0_70_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09101_ _09941_/A _09101_/B vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__or2_1
XANTENNA__08878__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07293_ _09767_/B _07293_/B vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ _09032_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_170_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12200__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12036__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold333 hold333/A vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold344 hold344/A vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold366 hold366/A vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold377 hold377/A vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11875__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout802 _12689_/S1 vssd1 vssd1 vccd1 vccd1 _12699_/S1 sky130_fd_sc_hd__clkbuf_8
Xhold388 hold388/A vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold399 hold399/A vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _13750_/A _13364_/B vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout813 _14489_/Q vssd1 vssd1 vccd1 vccd1 _12939_/S1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08168__C1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 _14488_/Q vssd1 vssd1 vccd1 vccd1 _12641_/S sky130_fd_sc_hd__buf_6
Xfanout835 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _12915_/S sky130_fd_sc_hd__buf_8
XFILLER_0_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12503__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 _13477_/A vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__buf_4
X_09865_ _10022_/B _10306_/A _09866_/C _09866_/D vssd1 vssd1 vccd1 vccd1 _09865_/X
+ sky130_fd_sc_hd__and4_1
Xfanout857 _13622_/C1 vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13375__B _13375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 _11681_/X vssd1 vssd1 vccd1 vccd1 _14484_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout868 _13487_/A vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout572_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08469__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _14218_/Q vssd1 vssd1 vccd1 vccd1 hold1011/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _06946_/Y vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__buf_6
XANTENNA__09380__A1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _13211_/X vssd1 vssd1 vccd1 vccd1 _15075_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _08816_/A _08816_/B _08816_/C vssd1 vssd1 vccd1 vccd1 _08820_/B sky130_fd_sc_hd__nand3_2
Xhold1033 _14618_/Q vssd1 vssd1 vccd1 vccd1 hold1033/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _10244_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09796_/Y sky130_fd_sc_hd__nor2_1
Xhold1044 _13505_/X vssd1 vssd1 vccd1 vccd1 _15263_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 _14008_/Q vssd1 vssd1 vccd1 vccd1 hold1055/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 _07526_/X vssd1 vssd1 vccd1 vccd1 _14151_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _14678_/Q vssd1 vssd1 vccd1 vccd1 hold1077/X sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _15145_/Q _09925_/A2 _08256_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _08747_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_90_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 _11925_/X vssd1 vssd1 vccd1 vccd1 _14746_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1099 _14660_/Q vssd1 vssd1 vccd1 vccd1 hold1099/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__A1 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_206 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13391__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_217 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12362__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ _08678_/A _08678_/B _08678_/C vssd1 vssd1 vccd1 vccd1 _08816_/A sky130_fd_sc_hd__and3_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11623__B _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ hold1707/X _13735_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07629_/X sky130_fd_sc_hd__mux2_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _11620_/A _11378_/D _10639_/C _10639_/D vssd1 vssd1 vccd1 vccd1 _10641_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08643__B1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _13586_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10751_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ _12294_/X _12326_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12310_/X sky130_fd_sc_hd__and3b_1
X_13290_ _13317_/A _13290_/B vssd1 vssd1 vccd1 vccd1 _15116_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12241_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_122_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_163_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ _14897_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11950__A0 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11123_ _15387_/Q _15290_/Q hold753/A _14391_/Q _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _11123_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_130_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07564__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ _11567_/A _15225_/Q _11055_/A vssd1 vssd1 vccd1 vccd1 _11054_/Y sky130_fd_sc_hd__nand3_1
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_178_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ _10005_/A _10005_/B vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__xnor2_2
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2290 _13469_/X vssd1 vssd1 vccd1 vccd1 _15228_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _14844_/CLK _14813_/D vssd1 vssd1 vccd1 vccd1 _14813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09123__A1 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_101_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13505__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09123__B2 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07134__A0 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14744_ _14926_/CLK _14744_/D vssd1 vssd1 vccd1 vccd1 _14744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08395__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _13711_/A1 hold773/X _11959_/S vssd1 vssd1 vccd1 vccd1 hold774/A sky130_fd_sc_hd__mux2_1
XANTENNA__09674__A2 _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06908__A _15345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07503__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ _11091_/B _10905_/X _10721_/X _10723_/Y vssd1 vssd1 vccd1 vccd1 _10907_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07685__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11887_ hold1267/X _13708_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 _11887_/X sky130_fd_sc_hd__mux2_1
X_14675_ _15062_/CLK hold446/X vssd1 vssd1 vccd1 vccd1 hold445/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10838_ _10840_/C vssd1 vssd1 vccd1 vccd1 _11015_/A sky130_fd_sc_hd__inv_2
X_13626_ input39/X _13634_/B vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_116_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12430__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ _08535_/B _09222_/B _13556_/X _13541_/A vssd1 vssd1 vccd1 vccd1 _13557_/X
+ sky130_fd_sc_hd__o211a_1
X_10769_ _11504_/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10769_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_137_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _15398_/Q _14533_/Q hold815/A _14757_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12508_/X sky130_fd_sc_hd__mux4_1
X_13488_ _13490_/A hold89/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__and2_1
XFILLER_0_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15227_ _15324_/CLK _15227_/D vssd1 vssd1 vccd1 vccd1 _15227_/Q sky130_fd_sc_hd__dfxtp_2
X_12439_ hold503/X hold1695/X hold1679/X hold1141/X _12460_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12439_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10419__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09954__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15158_ _15460_/CLK _15158_/D vssd1 vssd1 vccd1 vccd1 _15158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _14397_/CLK _14109_/D vssd1 vssd1 vccd1 vccd1 _14109_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13476__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15089_ _15089_/CLK hold308/X vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07980_ _07390_/A _07978_/Y _07979_/X _09925_/A2 _15136_/Q vssd1 vssd1 vccd1 vccd1
+ _07981_/C sky130_fd_sc_hd__a32o_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06931_ _14087_/Q vssd1 vssd1 vccd1 vccd1 _07875_/B sky130_fd_sc_hd__inv_2
XANTENNA__13195__B _13195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09650_ _10430_/B1 _09643_/Y _09645_/Y _09647_/Y _09649_/Y vssd1 vssd1 vccd1 vccd1
+ _09650_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_59_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08601_ _09008_/A _09860_/A _08470_/X _08383_/B _09858_/B vssd1 vssd1 vccd1 vccd1
+ _08607_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09581_ _10110_/A _10115_/A _09724_/C _09724_/D vssd1 vssd1 vccd1 vccd1 _09721_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_145_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12310__A_N _12294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12249__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08548__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _13384_/B vssd1 vssd1 vccd1 vccd1 _08532_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07676__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _08880_/A1 _08456_/Y _08458_/Y _08460_/Y _08462_/Y vssd1 vssd1 vccd1 vccd1
+ _08463_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_147_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ hold197/X _07475_/B vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__and2_1
XFILLER_0_147_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08394_ _08393_/A _08393_/B _08393_/C vssd1 vssd1 vccd1 vccd1 _08395_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07345_ _07345_/A _07345_/B _15327_/Q _15326_/Q vssd1 vssd1 vccd1 vccd1 _07362_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09848__B _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__A2 _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15429_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout418_A _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ _10827_/C _09726_/B vssd1 vssd1 vccd1 vccd1 _07277_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12274__B _13434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ _09013_/X _09015_/B vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_182_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10075__A _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09864__A _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A _14941_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13386__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout610 _15207_/Q vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__buf_6
Xfanout621 _10142_/A vssd1 vssd1 vccd1 vccd1 _09714_/A sky130_fd_sc_hd__buf_4
Xfanout632 _15201_/Q vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__clkbuf_8
X_09917_ _11288_/A1 _13395_/B _09807_/X vssd1 vssd1 vccd1 vccd1 _13448_/B sky130_fd_sc_hd__a21oi_4
Xfanout643 _15199_/Q vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__buf_4
XANTENNA__12488__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 _13715_/A1 vssd1 vssd1 vccd1 vccd1 _13748_/A1 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_97_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _14992_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout665 _15063_/Q vssd1 vssd1 vccd1 vccd1 hold2765/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout676 hold2728/X vssd1 vssd1 vccd1 vccd1 _13705_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__12583__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09848_ _10115_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__and2_1
Xfanout687 _15053_/Q vssd1 vssd1 vccd1 vccd1 _13700_/A1 sky130_fd_sc_hd__buf_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout698 _13727_/A1 vssd1 vssd1 vccd1 vccd1 _13661_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ _09780_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__and2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ hold1151/X _13664_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12335__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ hold475/A _14125_/Q _12791_/S vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__mux2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _13727_/A1 hold1983/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__mux2_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14460_ _15397_/CLK _14460_/D vssd1 vssd1 vccd1 vccd1 _14460_/Q sky130_fd_sc_hd__dfxtp_1
X_11672_ _13703_/A1 hold1565/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11672_/X sky130_fd_sc_hd__mux2_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ _11590_/A _11605_/B _10623_/C _10623_/D vssd1 vssd1 vccd1 vccd1 _10623_/Y
+ sky130_fd_sc_hd__nand4_4
X_13411_ _13459_/A _13411_/B vssd1 vssd1 vccd1 vccd1 _15199_/D sky130_fd_sc_hd__and2_1
XFILLER_0_154_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12412__A1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14391_ _15387_/CLK _14391_/D vssd1 vssd1 vccd1 vccd1 _14391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13060__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _14557_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13342_ _13342_/A _13342_/B vssd1 vssd1 vccd1 vccd1 _13343_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07559__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ _10553_/B _10553_/C _10553_/A vssd1 vssd1 vccd1 vccd1 _10554_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ input130/X fanout6/X fanout4/X input98/X vssd1 vssd1 vccd1 vccd1 _13273_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07278__B _14965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10485_ _11563_/A _11569_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _10652_/A
+ sky130_fd_sc_hd__nand4_2
X_15012_ _15177_/CLK _15012_/D vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
X_12224_ hold2710/X input1/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13172_/B sky130_fd_sc_hd__mux2_4
XANTENNA__09041__B1 _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13296__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _14984_/Q _12173_/A2 _12154_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12155_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07294__A _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _11645_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__nand2_1
X_12086_ _14983_/Q _12126_/B _12128_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12086_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_88_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15292_/CLK sky130_fd_sc_hd__clkbuf_16
X_11037_ _11037_/A _11037_/B _11037_/C vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12574__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A1 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11151__B2 _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13235__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ _06943_/A _12983_/X _12987_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12995_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _14791_/CLK hold968/X vssd1 vssd1 vccd1 vccd1 hold967/A sky130_fd_sc_hd__dfxtp_1
X_11939_ hold183/X hold2799/X _11943_/S vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__mux2_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ _15432_/CLK hold436/X vssd1 vssd1 vccd1 vccd1 hold435/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13609_ input61/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13609_/X sky130_fd_sc_hd__or2_1
XANTENNA__12403__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09804__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14589_ _15296_/CLK _14589_/D vssd1 vssd1 vccd1 vccd1 _14589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08572__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15423_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07130_ _13698_/A1 hold2231/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07130_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12954__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10965__A1 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__C _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10965__B2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07061_ _13666_/A1 hold1745/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07061_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput202 _14185_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[15] sky130_fd_sc_hd__buf_12
XFILLER_0_113_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12706__A2 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput213 _14195_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[25] sky130_fd_sc_hd__buf_12
XFILLER_0_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput224 _14176_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[6] sky130_fd_sc_hd__buf_12
XFILLER_0_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput235 _14440_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[16] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput246 _14450_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[26] sky130_fd_sc_hd__buf_12
Xoutput257 _14431_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[7] sky130_fd_sc_hd__buf_12
XFILLER_0_121_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput268 _14894_/Q vssd1 vssd1 vccd1 vccd1 out0[17] sky130_fd_sc_hd__buf_12
XFILLER_0_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10623__A _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput279 _14904_/Q vssd1 vssd1 vccd1 vccd1 out0[27] sky130_fd_sc_hd__buf_12
X_07963_ _07963_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__and2_1
XANTENNA__11438__B _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_79_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _14483_/CLK sky130_fd_sc_hd__clkbuf_16
X_09702_ _09701_/X _10010_/B _10110_/A _09702_/D vssd1 vssd1 vccd1 vccd1 _09704_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06914_ _06914_/A vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__inv_2
X_07894_ _07963_/A _07894_/B _07894_/C vssd1 vssd1 vccd1 vccd1 _07895_/A sky130_fd_sc_hd__and3_1
XANTENNA__11142__A1 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__B2 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ hold207/A _14318_/Q _14609_/Q _13978_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09633_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09850__C _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout368_A _07900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07992__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12317__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12269__B _13424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ _08516_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12642__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _09495_/A _13586_/B vssd1 vssd1 vccd1 vccd1 _09495_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout535_A _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08446_ hold229/A hold505/A _14599_/Q _13968_/Q _07816_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08446_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06982__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08377_ _08528_/D _08528_/B _09133_/A vssd1 vssd1 vccd1 vccd1 _08378_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_135_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07328_ _07328_/A _07328_/B _09205_/A _09619_/A vssd1 vssd1 vccd1 vccd1 _07328_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_163_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ _11614_/B _10108_/C vssd1 vssd1 vccd1 vccd1 _07261_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10270_ _11578_/A _14964_/Q _11573_/B _11580_/A vssd1 vssd1 vccd1 vccd1 _10293_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09574__A1 _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12224__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10184__A2 _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _07512_/Y vssd1 vssd1 vccd1 vccd1 _07544_/S sky130_fd_sc_hd__clkbuf_16
Xfanout451 _07981_/A vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__buf_4
Xfanout462 _12056_/S vssd1 vssd1 vccd1 vccd1 _12062_/S sky130_fd_sc_hd__clkbuf_8
Xfanout473 _13450_/A vssd1 vssd1 vccd1 vccd1 _13440_/S sky130_fd_sc_hd__buf_4
X_13960_ _15429_/CLK _13960_/D vssd1 vssd1 vccd1 vccd1 _13960_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout484 _11283_/S vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__clkbuf_16
Xfanout495 _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12644_/A1 sky130_fd_sc_hd__buf_8
X_12911_ _12917_/A1 _12910_/X _12950_/S0 vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07888__A1 _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ _15387_/CLK _13891_/D vssd1 vssd1 vccd1 vccd1 _13891_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12881__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12917_/A1 _12841_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07983__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12773_ hold239/A _14316_/Q hold541/A _13976_/Q _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12773_/X sky130_fd_sc_hd__mux4_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10644__B1 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14512_ _15444_/CLK hold550/X vssd1 vssd1 vccd1 vccd1 hold549/A sky130_fd_sc_hd__dfxtp_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ hold849/X _15064_/Q _11728_/S vssd1 vssd1 vccd1 vccd1 hold850/A sky130_fd_sc_hd__mux2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11655_ _13719_/A1 hold2251/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__mux2_1
X_14443_ _15313_/CLK _14443_/D vssd1 vssd1 vccd1 vccd1 _14443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07289__A _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10606_ _11578_/A _11577_/A _11573_/B _14966_/Q vssd1 vssd1 vccd1 vccd1 _10788_/A
+ sky130_fd_sc_hd__and4_1
X_11586_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14374_ _15440_/CLK _14374_/D vssd1 vssd1 vccd1 vccd1 _14374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13325_ input84/X fanout2/X _13324_/X vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__a21oi_1
X_10537_ _10362_/B _10364_/B _10534_/X _10535_/Y vssd1 vssd1 vccd1 vccd1 _10537_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13256_ input91/X fanout1/X _13255_/X vssd1 vssd1 vccd1 vccd1 _13257_/B sky130_fd_sc_hd__a21oi_1
X_10468_ _11586_/A _11614_/A _11623_/A vssd1 vssd1 vccd1 vccd1 _10468_/X sky130_fd_sc_hd__and3_1
XANTENNA__12244__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12207_ _12243_/A _12202_/X _12206_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _12208_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13187_ _13393_/A _13187_/B vssd1 vssd1 vccd1 vccd1 _15052_/D sky130_fd_sc_hd__and2_1
X_10399_ _10395_/Y _10397_/Y _10398_/X vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__a21o_2
XANTENNA__11372__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ _14880_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11973__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ hold2511/X _12099_/A2 _12068_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12069_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_1_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15394_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08525__C1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08540__A2 _12270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07471__B _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08300_ _08503_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__or2_1
XFILLER_0_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09280_ _09160_/A _09159_/B _09159_/A vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__08583__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08231_ _08230_/B _08230_/C _08230_/A vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ _08162_/A _08162_/B _08162_/C vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12483__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07113_ _14087_/Q _07114_/B vssd1 vssd1 vccd1 vccd1 _13502_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08093_ _08093_/A _08093_/B _08093_/C vssd1 vssd1 vccd1 vccd1 _08095_/B sky130_fd_sc_hd__or3_1
XFILLER_0_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08638__B1_N _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07044_ hold871/X _13748_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold872/A sky130_fd_sc_hd__mux2_1
XFILLER_0_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12235__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09100__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11168__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2801 _15051_/Q vssd1 vssd1 vccd1 vccd1 hold2801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2812 _12833_/X vssd1 vssd1 vccd1 vccd1 hold2812/X sky130_fd_sc_hd__dlygate4sd3_1
X_08995_ hold2739/X input7/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13187_/B sky130_fd_sc_hd__mux2_1
Xhold2823 _15051_/Q vssd1 vssd1 vccd1 vccd1 hold2823/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11883__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2834 _15301_/Q vssd1 vssd1 vccd1 vccd1 hold2834/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13104__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2845 _15349_/Q vssd1 vssd1 vccd1 vccd1 hold2845/X sky130_fd_sc_hd__dlygate4sd3_1
X_07946_ _07931_/Y _07936_/Y _07945_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _07947_/B sky130_fd_sc_hd__a221o_1
Xhold2856 _15315_/Q vssd1 vssd1 vccd1 vccd1 hold2856/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08758__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13383__B _13383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _07862_/C _14086_/Q _07875_/X _07876_/X vssd1 vssd1 vccd1 vccd1 _07878_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12863__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A _15197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08477__B _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09616_ _09616_/A _09616_/B vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08908__D _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09547_ _09547_/A _09547_/B _09547_/C vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__A1 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09478_ _09478_/A _09478_/B vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_136_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09492__B1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07601__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08429_ _08429_/A _08429_/B vssd1 vssd1 vccd1 vccd1 _08429_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10528__A _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11573_/A _11594_/B _11439_/C _11439_/D vssd1 vssd1 vccd1 vccd1 _11441_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08047__A1 _14428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11371_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13591__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ _10148_/A _10148_/C _10148_/B vssd1 vssd1 vccd1 vccd1 _10324_/C sky130_fd_sc_hd__a21bo_1
X_13110_ _13489_/A hold69/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__and2_1
X_14090_ _15293_/CLK _14090_/D vssd1 vssd1 vccd1 vccd1 _14090_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_15_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13558__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ hold629/A hold797/A _13041_/S vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__mux2_1
X_10253_ _15414_/Q _14549_/Q _14709_/Q _14773_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10253_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09642__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _11351_/B _10830_/B _10356_/C _10183_/A vssd1 vssd1 vccd1 vccd1 _10185_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11793__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14992_ _14992_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 _14992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07572__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13943_ _15056_/CLK _13943_/D vssd1 vssd1 vccd1 vccd1 _13943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12854__A1 _13395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07291__B _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ _14569_/CLK _13874_/D vssd1 vssd1 vccd1 vccd1 _13874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12606__A1 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ _12821_/X _12822_/X _12824_/X _12823_/X _12844_/A1 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12826_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13513__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08286__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09483__B1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _13106_/A1 _13157_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12757_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_189_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ hold1375/X _13661_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11707_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12687_ _12689_/S1 _12684_/X _12686_/X vssd1 vssd1 vccd1 vccd1 _12687_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14426_ _15304_/CLK _14426_/D vssd1 vssd1 vccd1 vccd1 _14426_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_86_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11638_ _11469_/Y _11473_/C _11637_/Y vssd1 vssd1 vccd1 vccd1 _11638_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13031__A1 _07355_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11968__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13749__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14357_ _15385_/CLK hold736/X vssd1 vssd1 vccd1 vccd1 hold735/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ _11569_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nand2_1
Xhold707 hold707/A vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ _13317_/A _13308_/B vssd1 vssd1 vccd1 vccd1 _15122_/D sky130_fd_sc_hd__nor2_1
Xhold718 hold718/A vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13468__B _13468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold729 hold729/A vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ _14651_/CLK hold594/X vssd1 vssd1 vccd1 vccd1 hold593/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10173__A _14942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ _15353_/Q _15352_/Q _13239_/C _13239_/D vssd1 vssd1 vccd1 vccd1 _13241_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09633__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__B1 _14490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2108 _11717_/X vssd1 vssd1 vccd1 vccd1 _14513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2119 _14380_/Q vssd1 vssd1 vccd1 vccd1 hold2119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07800_ hold1127/X _13738_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 _07800_/X sky130_fd_sc_hd__mux2_1
X_08780_ _08901_/A _08892_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _08780_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1407 _14732_/Q vssd1 vssd1 vccd1 vccd1 hold1407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1418 _13511_/X vssd1 vssd1 vccd1 vccd1 _15269_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 _14296_/Q vssd1 vssd1 vccd1 vccd1 hold1429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07731_ hold407/X _13671_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold408/A sky130_fd_sc_hd__mux2_1
XFILLER_0_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09710__A1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07662_ hold1265/X hold169/X _07676_/S vssd1 vssd1 vccd1 vccd1 _07662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_189_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09401_ _10129_/A _10022_/A _09247_/X _09248_/X _10126_/A vssd1 vssd1 vccd1 vccd1
+ _09406_/A sky130_fd_sc_hd__a32o_1
XANTENNA__12506__A1_N _08253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07593_ _13732_/A1 hold1467/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07593_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _09195_/Y _09197_/Y _09330_/Y _09331_/X vssd1 vssd1 vccd1 vccd1 _09335_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13270__A1 input160/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09263_ _09449_/A vssd1 vssd1 vccd1 vccd1 _09264_/D sky130_fd_sc_hd__inv_2
XFILLER_0_168_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08214_ _08214_/A _08297_/B _08214_/C vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__and3_1
XFILLER_0_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ _09328_/A _09194_/B vssd1 vssd1 vccd1 vccd1 _09196_/B sky130_fd_sc_hd__and2_1
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09226__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11878__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08145_ _08144_/B _08144_/C _08144_/A vssd1 vssd1 vccd1 vccd1 _08147_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08124__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout400_A _07577_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12781__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ _08075_/B _10507_/A _11550_/A _08892_/A vssd1 vssd1 vccd1 vccd1 _08077_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13378__B _13378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__B _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07027_ hold1569/X _13665_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07027_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13394__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2620 _08262_/X vssd1 vssd1 vccd1 vccd1 _14431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2631 _09632_/X vssd1 vssd1 vccd1 vccd1 _14443_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2642 _14444_/Q vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08978_ _08981_/A _08975_/X _08977_/X vssd1 vssd1 vccd1 vccd1 _08978_/Y sky130_fd_sc_hd__o21ai_1
Xhold2653 _14979_/Q vssd1 vssd1 vccd1 vccd1 hold2653/X sky130_fd_sc_hd__buf_2
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2664 _09223_/X vssd1 vssd1 vccd1 vccd1 _14440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2675 _12030_/X vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1930 _07522_/X vssd1 vssd1 vccd1 vccd1 _14147_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2686 _14822_/Q vssd1 vssd1 vccd1 vccd1 hold2686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _13865_/Q hold681/A _13833_/Q _13801_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07929_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12836__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1941 _13913_/Q vssd1 vssd1 vccd1 vccd1 hold1941/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2697 _12062_/X vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1952 _11915_/X vssd1 vssd1 vccd1 vccd1 _14736_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1963 _14383_/Q vssd1 vssd1 vccd1 vccd1 hold1963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1974 _07407_/X vssd1 vssd1 vccd1 vccd1 _14037_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ hold599/A hold835/A hold493/A hold999/A _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _10941_/B sky130_fd_sc_hd__mux4_1
Xhold1985 _14369_/Q vssd1 vssd1 vccd1 vccd1 hold1985/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08060__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1996 _07676_/X vssd1 vssd1 vccd1 vccd1 _14297_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10942__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ _10686_/B _10688_/B _10686_/A vssd1 vssd1 vccd1 vccd1 _10872_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ hold997/A _13938_/Q _12735_/S vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08268__A1 _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13261__A1 input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13590_ _13590_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13590_/X sky130_fd_sc_hd__or2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11498__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ hold499/A _14243_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13549__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _15389_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold707/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13013__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12447__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ _14787_/Q _14499_/Q hold995/A _14723_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12472_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14211_ _15045_/CLK hold578/X vssd1 vssd1 vccd1 vccd1 hold577/A sky130_fd_sc_hd__dfxtp_1
X_11423_ _11420_/X _11421_/Y _11177_/B _11179_/B vssd1 vssd1 vccd1 vccd1 _11449_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15191_ _15191_/CLK _15191_/D vssd1 vssd1 vccd1 vccd1 _15191_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12998__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _11354_/A _11354_/B _11354_/C vssd1 vssd1 vccd1 vccd1 _11518_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07567__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _15397_/CLK hold752/X vssd1 vssd1 vccd1 vccd1 hold751/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10305_ _11564_/A _11606_/A _10306_/C _10306_/D vssd1 vssd1 vccd1 vccd1 _10305_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_123_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07286__B _14972_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14073_ _15356_/CLK _14073_/D vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
X_11285_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13024_ _13890_/Q hold293/A _13858_/Q _13826_/Q _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _13024_/X sky130_fd_sc_hd__mux4_1
X_10236_ _13749_/A _13452_/B _10235_/X vssd1 vssd1 vccd1 vccd1 _10236_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13508__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _11335_/A _10338_/D _10165_/Y _10343_/A vssd1 vssd1 vccd1 vccd1 _10169_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07506__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11536__B _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10098_ _11504_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10098_/Y sky130_fd_sc_hd__nor2_1
X_14975_ _14975_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 _14975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07929__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ _15427_/CLK _13926_/D vssd1 vssd1 vccd1 vccd1 _13926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08051__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10933__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ _15454_/CLK _13857_/D vssd1 vssd1 vccd1 vccd1 _13857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12808_ hold1719/X _14545_/Q hold933/A hold1173/X _12841_/S _06942_/A vssd1 vssd1
+ vccd1 vccd1 _12808_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08259__A1 _14430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13252__A1 input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13788_ _06907_/A _13792_/A2 _11685_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _15346_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12739_ _14283_/Q hold1203/X hold2805/X hold873/X _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12739_/X sky130_fd_sc_hd__mux4_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12086__C _12128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13004__A1 _10918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15458_ _15458_/CLK hold362/X vssd1 vssd1 vccd1 vccd1 hold361/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11698__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ _14409_/CLK hold748/X vssd1 vssd1 vccd1 vccd1 hold747/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13555__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12989__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15389_ _15389_/CLK hold368/X vssd1 vssd1 vccd1 vccd1 hold367/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold504 hold504/A vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 hold515/A vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13198__B _13198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__B2 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold526 hold526/A vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 hold537/A vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 hold548/A vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09950_ _15412_/Q _14547_/Q hold491/A _14771_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _09950_/X sky130_fd_sc_hd__mux4_1
Xhold559 hold559/A vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11318__A1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08901_ _08901_/A _09726_/B _08901_/C vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09881_ _09881_/A _09881_/B _09881_/C vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__and3_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08829_/Y _08830_/X _08721_/B _08721_/Y vssd1 vssd1 vccd1 vccd1 _08833_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _07595_/X vssd1 vssd1 vccd1 vccd1 _14219_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 _14690_/Q vssd1 vssd1 vccd1 vccd1 hold1215/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _11719_/X vssd1 vssd1 vccd1 vccd1 _14515_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1237 _13817_/Q vssd1 vssd1 vccd1 vccd1 hold1237/X sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ _14279_/Q _14215_/Q _14151_/Q _14469_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08764_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12818__A1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1248 _11845_/X vssd1 vssd1 vccd1 vccd1 _14668_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 _15084_/Q vssd1 vssd1 vccd1 vccd1 hold1259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07714_ hold595/X _13687_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold596/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ _08694_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _08697_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07940__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10777__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ hold619/X _12329_/A _07660_/S vssd1 vssd1 vccd1 vccd1 hold620/A sky130_fd_sc_hd__mux2_1
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout448_A _07389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13243__A1 input129/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _13404_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _14201_/D sky130_fd_sc_hd__and2_1
XFILLER_0_211_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07151__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12277__B _12277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09315_ _09314_/B _09314_/C _09314_/A vssd1 vssd1 vccd1 vccd1 _09317_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout615_A _15206_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09246_ _10129_/A _10022_/A vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06990__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08771__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13389__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _09178_/A _09178_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__and3_1
XFILLER_0_161_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14923__D _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08958__C1 _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ _14659_/Q _13932_/Q _15433_/Q _13900_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08129_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _08760_/A _08059_/B vssd1 vssd1 vccd1 vccd1 _08059_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12506__B1 _13147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _10885_/B _10887_/B _11067_/X _11068_/Y vssd1 vssd1 vccd1 vccd1 _11070_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput102 in1[14] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__clkbuf_1
X_10021_ _10022_/B _10304_/C _10304_/D _10022_/A vssd1 vssd1 vccd1 vccd1 _10024_/B
+ sky130_fd_sc_hd__a22oi_2
Xinput113 in1[24] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12232__S _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput124 in1[5] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08281__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput135 in2[15] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__clkbuf_2
Xinput146 in2[25] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__clkbuf_2
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2450 hold2842/X vssd1 vssd1 vccd1 vccd1 _07428_/A sky130_fd_sc_hd__buf_1
Xinput157 in2[6] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__clkbuf_2
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2461 _14870_/Q vssd1 vssd1 vccd1 vccd1 hold2461/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09107__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2472 _12165_/X vssd1 vssd1 vccd1 vccd1 _14893_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2483 _14875_/Q vssd1 vssd1 vccd1 vccd1 hold2483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2494 _12119_/X vssd1 vssd1 vccd1 vccd1 _14871_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1760 _06979_/X vssd1 vssd1 vccd1 vccd1 _13798_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1771 _14510_/Q vssd1 vssd1 vccd1 vccd1 hold1771/X sky130_fd_sc_hd__dlygate4sd3_1
X_14760_ _15042_/CLK _14760_/D vssd1 vssd1 vccd1 vccd1 _14760_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ hold1583/X _13661_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11972_/X sky130_fd_sc_hd__mux2_1
Xhold1782 _07772_/X vssd1 vssd1 vccd1 vccd1 _14388_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1793 _13911_/Q vssd1 vssd1 vccd1 vccd1 hold1793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_2_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ hold1659/X _13711_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13711_/X sky130_fd_sc_hd__mux2_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _11108_/D _10923_/B vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__xnor2_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _15394_/CLK _14691_/D vssd1 vssd1 vccd1 vccd1 _14691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13642_ input53/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13642_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10854_ _10663_/X _10668_/A _10852_/X _10853_/Y vssd1 vssd1 vccd1 vccd1 _10856_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13234__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07061__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _06916_/A _13586_/B _13572_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13573_/X
+ sky130_fd_sc_hd__o211a_1
X_10785_ _11573_/B _10784_/X _10783_/X vssd1 vssd1 vccd1 vccd1 _10787_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08110__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15312_ _15316_/CLK _15312_/D vssd1 vssd1 vccd1 vccd1 _15312_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _13870_/Q hold421/A hold905/A _13806_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12524_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13299__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15243_ _15243_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
X_12455_ _12327_/A hold2730/X _12452_/X vssd1 vssd1 vccd1 vccd1 _13145_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_48_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07297__A _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ _11168_/A _11606_/B _11570_/B _11407_/A vssd1 vssd1 vccd1 vccd1 _11408_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15174_ _15177_/CLK _15174_/D vssd1 vssd1 vccd1 vccd1 _15174_/Q sky130_fd_sc_hd__dfxtp_2
X_12386_ _12642_/A1 _12385_/X _12644_/A1 vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ _14612_/CLK _14125_/D vssd1 vssd1 vccd1 vccd1 _14125_/Q sky130_fd_sc_hd__dfxtp_1
X_11337_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14056_ _15351_/CLK _14056_/D vssd1 vssd1 vccd1 vccd1 _14056_/Q sky130_fd_sc_hd__dfxtp_1
X_11268_ _11039_/Y _11081_/B _11080_/A vssd1 vssd1 vccd1 vccd1 _11269_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09913__A1 _11474_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13007_ _13171_/A _13007_/B vssd1 vssd1 vccd1 vccd1 _14968_/D sky130_fd_sc_hd__nor2_1
X_10219_ _10266_/B _10220_/B _10220_/C vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11199_ _11197_/X _11199_/B vssd1 vssd1 vccd1 vccd1 _11200_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11981__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14958_ _14958_/CLK _14958_/D vssd1 vssd1 vccd1 vccd1 _14958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _15442_/CLK _13909_/D vssd1 vssd1 vccd1 vccd1 _13909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10597__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889_ _14889_/CLK _14889_/D vssd1 vssd1 vccd1 vccd1 _14889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07430_ _07430_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14060_/D sky130_fd_sc_hd__and2_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09429__B1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07361_ _13468_/A _07360_/Y _14022_/Q vssd1 vssd1 vccd1 vccd1 _07846_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09100_ _14797_/Q _14509_/Q _14637_/Q _14733_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09101_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13701__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07292_ _11542_/B _10115_/D vssd1 vssd1 vccd1 vccd1 _07293_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09031_ _09030_/A _09030_/B _09030_/C vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2747_A _15181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07919__B _07919_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__B1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13002__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__A1 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__B2 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold334 hold334/A vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold345 hold345/A vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 hold367/A vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 hold378/A vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold389 hold389/A vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _13364_/B sky130_fd_sc_hd__or2_1
Xfanout803 _12689_/S1 vssd1 vssd1 vccd1 vccd1 _12674_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout814 _14489_/Q vssd1 vssd1 vccd1 vccd1 _13074_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout825 _12365_/S0 vssd1 vssd1 vccd1 vccd1 _12466_/S sky130_fd_sc_hd__buf_6
XANTENNA__09365__C1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A _07610_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout836 _13066_/S vssd1 vssd1 vccd1 vccd1 _12866_/S sky130_fd_sc_hd__buf_6
XANTENNA__12052__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ _09864_/A _10022_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _09866_/D
+ sky130_fd_sc_hd__nand4_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 _13481_/A vssd1 vssd1 vccd1 vccd1 _13386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout858 _13622_/C1 vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__buf_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _13827_/Q vssd1 vssd1 vccd1 vccd1 hold1001/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _13492_/A vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__buf_4
Xhold1012 _07594_/X vssd1 vssd1 vccd1 vccd1 _14218_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07146__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__A2 _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ _08814_/B _08814_/C _08814_/A vssd1 vssd1 vccd1 vccd1 _08816_/C sky130_fd_sc_hd__a21o_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _15364_/Q vssd1 vssd1 vccd1 vccd1 hold1023/X sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ hold383/A _14255_/Q _14415_/Q _14127_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09796_/B sky130_fd_sc_hd__mux4_1
Xhold1034 _11793_/X vssd1 vssd1 vccd1 vccd1 _14618_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout565_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 _13884_/Q vssd1 vssd1 vccd1 vccd1 hold1045/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _07201_/X vssd1 vssd1 vccd1 vccd1 _14008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 _14543_/Q vssd1 vssd1 vccd1 vccd1 hold1067/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06985__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08746_ _08746_/A _08746_/B vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__xnor2_1
Xhold1078 _11855_/X vssd1 vssd1 vccd1 vccd1 _14678_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08766__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 _13840_/Q vssd1 vssd1 vccd1 vccd1 hold1089/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13391__B _13391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_218 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08677_/A _08893_/A _09866_/B _09864_/C vssd1 vssd1 vccd1 vccd1 _08678_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA_fanout732_A _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12288__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07628_ hold1061/X _13734_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07628_/X sky130_fd_sc_hd__mux2_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08891__A1 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08891__B2 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09515__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07559_ _13393_/A hold143/X vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _10746_/B _10570_/B vssd1 vssd1 vccd1 vccd1 _13367_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ _14798_/Q _14510_/Q hold351/A _14734_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09230_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13075__S0 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12240_ _12247_/A _12235_/X _12239_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _12241_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ hold2593/X _12173_/A2 _12170_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12171_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12751__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _11507_/A _11119_/X _11121_/X vssd1 vssd1 vccd1 vccd1 _11122_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13566__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold890 hold890/A vssd1 vssd1 vccd1 vccd1 hold890/X sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ _11567_/A _15225_/Q vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__nand2_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10271__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _10005_/A _10005_/B vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__and2_1
XANTENNA__07056__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2280 _07106_/X vssd1 vssd1 vccd1 vccd1 _13919_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2291 _13964_/Q vssd1 vssd1 vccd1 vccd1 hold2291/X sky130_fd_sc_hd__dlygate4sd3_1
X_14812_ _15389_/CLK hold370/X vssd1 vssd1 vccd1 vccd1 hold369/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08676__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12889__S0 _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09123__A2 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1590 _11778_/X vssd1 vssd1 vccd1 vccd1 _14603_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14743_ _14791_/CLK _14743_/D vssd1 vssd1 vccd1 vccd1 _14743_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12663__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _13743_/A1 hold2035/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__mux2_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08395__B _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10906_ _10721_/X _10723_/Y _11091_/B _10905_/X vssd1 vssd1 vccd1 vccd1 _11098_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_156_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14674_ _15090_/CLK hold922/X vssd1 vssd1 vccd1 vccd1 hold921/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ hold325/X _15060_/Q _11893_/S vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ input38/X _13625_/B _13625_/C vssd1 vssd1 vccd1 vccd1 _15340_/D sky130_fd_sc_hd__and3_1
XFILLER_0_13_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10837_ _11605_/A _11570_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _10840_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12926__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13521__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08634__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ _14434_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13556_/X sky130_fd_sc_hd__or2_1
XANTENNA__06924__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _14293_/Q _14229_/Q hold633/A _14483_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10769_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09300__A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__A1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _12607_/A _12507_/B vssd1 vssd1 vccd1 vccd1 _14948_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ _13487_/A hold9/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__and2_1
XFILLER_0_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10699_ _11561_/A _11542_/B _11564_/B _14947_/Q vssd1 vssd1 vccd1 vccd1 _10700_/D
+ sky130_fd_sc_hd__a22o_1
X_15226_ _15226_/CLK _15226_/D vssd1 vssd1 vccd1 vccd1 _15226_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12438_ _12642_/B1 _12433_/X _12437_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12445_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11976__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15157_ _15423_/CLK _15157_/D vssd1 vssd1 vccd1 vccd1 _15157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12369_ _13864_/Q _13992_/Q _12566_/S vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ _15392_/CLK hold518/X vssd1 vssd1 vccd1 vccd1 hold517/A sky130_fd_sc_hd__dfxtp_1
X_15088_ _15377_/CLK _15088_/D vssd1 vssd1 vccd1 vccd1 _15088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07474__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14039_ _15229_/CLK _14039_/D vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
X_06930_ _14086_/Q vssd1 vssd1 vccd1 vccd1 _07875_/C sky130_fd_sc_hd__inv_2
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08608_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09580_ _10115_/A _09724_/C _09724_/D _10110_/A vssd1 vssd1 vccd1 vccd1 _09584_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08531_ _12258_/S _08569_/C _08530_/Y _08525_/X hold2589/X vssd1 vssd1 vccd1 vccd1
+ _13384_/B sky130_fd_sc_hd__o311a_4
XANTENNA__08548__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08462_ _12243_/A _08461_/X _08880_/A1 vssd1 vssd1 vccd1 vccd1 _08462_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ _13535_/B hold105/X vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__and2_1
X_08393_ _08393_/A _08393_/B _08393_/C vssd1 vssd1 vccd1 vccd1 _08395_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07344_ _06920_/A _07343_/X _07342_/X vssd1 vssd1 vccd1 vccd1 _07344_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_190_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07275_ _10827_/C _09726_/B vssd1 vssd1 vccd1 vccd1 _09075_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10432__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09014_ _09011_/Y _09012_/X _08892_/X _08894_/X vssd1 vssd1 vccd1 vccd1 _09015_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12185__A1 hold2535/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11886__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09864__B _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13386__B _13386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12290__B _13466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout682_A _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _15211_/Q vssd1 vssd1 vccd1 vccd1 _09676_/D sky130_fd_sc_hd__clkbuf_8
Xfanout611 _09708_/B vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__buf_6
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09916_ _11287_/S _09914_/Y _09915_/X _09913_/X vssd1 vssd1 vccd1 vccd1 _13395_/B
+ sky130_fd_sc_hd__a31o_4
Xfanout622 _10142_/A vssd1 vssd1 vccd1 vccd1 _11573_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout633 _15201_/Q vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__buf_2
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09889__B1 _09888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout644 _10002_/C vssd1 vssd1 vccd1 vccd1 _11577_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout655 _15068_/Q vssd1 vssd1 vccd1 vccd1 _13715_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__09353__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 _13742_/A1 vssd1 vssd1 vccd1 vccd1 _11921_/A0 sky130_fd_sc_hd__clkbuf_4
X_09847_ _09847_/A _10005_/A vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__or2_1
Xfanout677 _13704_/A1 vssd1 vssd1 vccd1 vccd1 _13671_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 _13732_/A1 vssd1 vssd1 vccd1 vccd1 _13666_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout699 hold183/X vssd1 vssd1 vccd1 vccd1 _13727_/A1 sky130_fd_sc_hd__buf_4
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12510__S _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09778_/A _09930_/A vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__xnor2_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07604__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08729_ _08621_/Y _08623_/Y _08727_/Y _08728_/X vssd1 vssd1 vccd1 vccd1 _08841_/A
+ sky130_fd_sc_hd__o211ai_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _13693_/A1 hold749/X _11745_/S vssd1 vssd1 vccd1 vccd1 hold750/A sky130_fd_sc_hd__mux2_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11671_ _13735_/A1 hold587/X _11684_/S vssd1 vssd1 vccd1 vccd1 hold588/A sky130_fd_sc_hd__mux2_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13410_ _07919_/A _12262_/B _13468_/A vssd1 vssd1 vccd1 vccd1 _13411_/B sky130_fd_sc_hd__mux2_1
X_10622_ _11598_/A _11569_/B _11563_/B _11597_/A vssd1 vssd1 vccd1 vccd1 _10623_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14390_ _15289_/CLK _14390_/D vssd1 vssd1 vccd1 vccd1 _14390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ _13369_/A _13341_/B vssd1 vssd1 vccd1 vccd1 _15133_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10553_ _10553_/A _10553_/B _10553_/C vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__or3_1
XFILLER_0_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13048__S0 _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13272_ _13287_/A _13272_/B vssd1 vssd1 vccd1 vccd1 _15110_/D sky130_fd_sc_hd__nor2_1
X_10484_ _10285_/B _10287_/B _10285_/A vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _15268_/CLK _15011_/D vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__dfxtp_1
X_12223_ _13374_/B vssd1 vssd1 vccd1 vccd1 _12223_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09041__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _12154_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__or2_1
XFILLER_0_159_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11105_ _11645_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__or2_1
XANTENNA__07294__B _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12479__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13676__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ hold2469/X _12099_/A2 _12084_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12085_/X
+ sky130_fd_sc_hd__o211a_1
X_11036_ _11037_/A _11037_/B _11037_/C vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08001__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11151__A2 _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13516__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _13024_/S1 _12984_/X _12986_/X vssd1 vssd1 vccd1 vccd1 _12987_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08304__B1 _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14726_ _15270_/CLK _14726_/D vssd1 vssd1 vccd1 vccd1 _14726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11938_ _13693_/A1 hold1521/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11938_/X sky130_fd_sc_hd__mux2_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14657_ _14754_/CLK _14657_/D vssd1 vssd1 vccd1 vccd1 _14657_/Q sky130_fd_sc_hd__dfxtp_1
X_11869_ hold1289/X _13657_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_157_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13608_ _06913_/A _13625_/C _13607_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14588_ _15292_/CLK hold228/X vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12403__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13539_ _07908_/A _13797_/A2 _13538_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _13539_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13039__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10965__A2 _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08291__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07060_ _13665_/A1 hold1859/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07060_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12167__A1 hold2439/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15209_ _15226_/CLK _15209_/D vssd1 vssd1 vccd1 vccd1 _15209_/Q sky130_fd_sc_hd__dfxtp_4
Xoutput203 _14186_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[16] sky130_fd_sc_hd__buf_12
XANTENNA__13487__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput214 _14196_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[26] sky130_fd_sc_hd__buf_12
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput225 _14177_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[7] sky130_fd_sc_hd__buf_12
XFILLER_0_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput236 _14441_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[17] sky130_fd_sc_hd__buf_12
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput247 _14451_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[27] sky130_fd_sc_hd__buf_12
XANTENNA__09583__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput258 _14432_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[8] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput269 _14895_/Q vssd1 vssd1 vccd1 vccd1 out0[18] sky130_fd_sc_hd__buf_12
XANTENNA__10623__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07962_ _07963_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11438__C _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _09846_/B _10002_/C _10283_/C _10115_/D vssd1 vssd1 vccd1 vccd1 _09701_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__11678__A0 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ _06913_/A vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__inv_2
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07893_ _07963_/A _07894_/B _07894_/C vssd1 vssd1 vccd1 vccd1 _07893_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11142__A2 _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _09498_/A _13586_/B _09631_/Y _13579_/C1 vssd1 vssd1 vccd1 vccd1 _09632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07897__A2 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09850__D _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _10115_/D _09427_/B _09562_/X vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_167_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08514_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08516_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_162_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10102__B1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _09494_/A1 _09357_/Y _09493_/X vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10653__A1 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10653__B2 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ _08545_/B _08444_/Y _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08541_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout430_A _11796_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout528_A _15425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ _13512_/A0 _12260_/A2 _12259_/A1 _13181_/B _08374_/Y vssd1 vssd1 vccd1 vccd1
+ _08376_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_190_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12285__B _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07327_ _10600_/A _07327_/B _07951_/A vssd1 vssd1 vccd1 vccd1 _07329_/C sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_177_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_57_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ _08846_/B _07258_/B vssd1 vssd1 vccd1 vccd1 _07320_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_131_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13397__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14931__D _14931_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ hold1887/X _13657_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07189_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08457__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11118__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _11796_/Y vssd1 vssd1 vccd1 vccd1 _11828_/S sky130_fd_sc_hd__clkbuf_16
Xfanout441 _08441_/B vssd1 vssd1 vccd1 vccd1 _09222_/B sky130_fd_sc_hd__buf_4
Xfanout452 _13636_/B vssd1 vssd1 vccd1 vccd1 _13634_/B sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_115_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _07045_/X vssd1 vssd1 vccd1 vccd1 _07061_/S sky130_fd_sc_hd__clkbuf_16
Xfanout474 _13466_/A vssd1 vssd1 vccd1 vccd1 _13450_/A sky130_fd_sc_hd__buf_4
Xfanout485 _07854_/Y vssd1 vssd1 vccd1 vccd1 _08526_/B sky130_fd_sc_hd__buf_8
X_12910_ hold771/A _13950_/Q _12915_/S vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__mux2_1
Xfanout496 _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12700_/S0 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07888__A2 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ _14483_/CLK _13890_/D vssd1 vssd1 vccd1 vccd1 _13890_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12881__A2 _13162_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12841_ hold383/A _14255_/Q _12841_/S vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__mux2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12772_ _14799_/Q _14511_/Q _14639_/Q _14735_/Q _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12772_/X sky130_fd_sc_hd__mux4_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14511_ _15376_/CLK _14511_/D vssd1 vssd1 vccd1 vccd1 _14511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10644__A1 _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ hold683/X hold2765/A _11728_/S vssd1 vssd1 vccd1 vccd1 hold684/A sky130_fd_sc_hd__mux2_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__B2 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12476__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11380__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _15313_/CLK _14442_/D vssd1 vssd1 vccd1 vccd1 _14442_/Q sky130_fd_sc_hd__dfxtp_1
X_11654_ _13718_/A1 hold2173/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11654_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10605_ _11577_/A _11573_/B _14966_/Q _11578_/A vssd1 vssd1 vccd1 vccd1 _10605_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07289__B _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14373_ _15080_/CLK _14373_/D vssd1 vssd1 vccd1 vccd1 _14373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11585_ _11381_/A _11381_/B _11379_/B vssd1 vssd1 vccd1 vccd1 _11587_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ input148/X fanout5/X fanout3/X input116/X vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__a22o_1
X_10536_ _10362_/B _10364_/B _10534_/X _10535_/Y vssd1 vssd1 vccd1 vccd1 _10536_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_134_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output182_A _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12149__A1 hold2602/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13255_ input155/X fanout6/X fanout4/X input123/X vssd1 vssd1 vccd1 vccd1 _13255_/X
+ sky130_fd_sc_hd__a22o_1
X_10467_ _10467_/A _10635_/A _10467_/C vssd1 vssd1 vccd1 vccd1 _10502_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_126_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12415__S _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12244__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07509__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _12231_/A _12203_/X _12205_/X vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__a21o_1
X_13186_ _13481_/A _13186_/B vssd1 vssd1 vccd1 vccd1 _15051_/D sky130_fd_sc_hd__and2_1
X_10398_ _12221_/B _10261_/Y _10262_/X _11474_/A2 hold2792/X vssd1 vssd1 vccd1 vccd1
+ _10398_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_209_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11372__A2 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ hold2548/X _12195_/A2 _12136_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12137_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13649__A1 _07448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09948__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12068_ _12068_/A _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12068_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_205_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11019_ _11018_/B _11201_/A _09075_/A vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_189_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14709_ _15408_/CLK _14709_/D vssd1 vssd1 vccd1 vccd1 _14709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08583__B _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _08230_/A _08230_/B _08230_/C vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__and3_1
XFILLER_0_129_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12388__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2562_A _14987_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08162_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_173_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12483__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ _13748_/A1 hold2003/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07112_/X sky130_fd_sc_hd__mux2_1
X_08092_ _08093_/A _08093_/B _08093_/C vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07043_ hold2045/X _13681_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 _07043_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09005__A1 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12235__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09100__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2802 _14208_/Q vssd1 vssd1 vccd1 vccd1 hold2802/X sky130_fd_sc_hd__dlygate4sd3_1
X_08994_ _11320_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _08994_/Y sky130_fd_sc_hd__nor2_1
Xhold2813 _14527_/Q vssd1 vssd1 vccd1 vccd1 hold2813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2824 _15333_/Q vssd1 vssd1 vccd1 vccd1 hold2824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2835 _15335_/Q vssd1 vssd1 vccd1 vccd1 hold2835/X sky130_fd_sc_hd__dlygate4sd3_1
X_07945_ _08564_/A1 _07938_/Y _07940_/Y _07942_/Y _07944_/Y vssd1 vssd1 vccd1 vccd1
+ _07945_/X sky130_fd_sc_hd__o32a_1
XANTENNA__09939__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2846 _15305_/Q vssd1 vssd1 vccd1 vccd1 hold2846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2857 _15348_/Q vssd1 vssd1 vccd1 vccd1 hold2857/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11115__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _07355_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12060__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ _15341_/Q _07875_/C _14090_/Q _06908_/Y vssd1 vssd1 vccd1 vccd1 _07876_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07154__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _09760_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09616_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_211_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout645_A _15199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09546_ _09673_/B _09545_/C _09545_/A vssd1 vssd1 vccd1 vccd1 _09547_/C sky130_fd_sc_hd__a21o_1
XANTENNA__06993__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09477_ _09762_/A _09762_/B _09762_/C _09476_/X vssd1 vssd1 vccd1 vccd1 _09478_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08295__A2 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout812_A _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ _08428_/A _08428_/B vssd1 vssd1 vccd1 vccd1 _08429_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10528__B _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09244__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ hold339/A _15270_/Q hold889/A _14371_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08359_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_163_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _11370_/A _11370_/B vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ _10320_/B _10320_/C _10320_/A vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12000__A0 _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ hold489/X hold1239/X _13091_/S vssd1 vssd1 vccd1 vccd1 _13040_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10252_ _10252_/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10252_/Y sky130_fd_sc_hd__nor2_1
X_10183_ _10183_/A _11351_/B _10830_/B _10356_/C vssd1 vssd1 vccd1 vccd1 _10185_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_100_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13574__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _15247_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 _14991_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13066__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11375__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13942_ _15377_/CLK _13942_/D vssd1 vssd1 vccd1 vccd1 _13942_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12854__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07064__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08387__C _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13873_ _15080_/CLK _13873_/D vssd1 vssd1 vccd1 vccd1 _13873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12824_ _13882_/Q hold617/A hold659/A _13818_/Q _12915_/S _12939_/S1 vssd1 vssd1
+ vccd1 vccd1 _12824_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12606__A2 _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12755_ _13080_/A1 _12754_/X _12752_/X vssd1 vssd1 vccd1 vccd1 _13157_/B sky130_fd_sc_hd__a21oi_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09483__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ hold2099/X _13512_/A0 _11712_/S vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12686_ _12692_/A1 _12685_/X _12700_/S0 vssd1 vssd1 vccd1 vccd1 _12686_/X sky130_fd_sc_hd__a21o_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14425_ _15456_/CLK hold886/X vssd1 vssd1 vccd1 vccd1 hold885/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11637_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14356_ _14971_/CLK _14356_/D vssd1 vssd1 vccd1 vccd1 _14356_/Q sky130_fd_sc_hd__dfxtp_1
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13749__B _13749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07797__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13307_ input78/X fanout2/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13308_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold708 hold708/A vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ _10519_/A _10519_/B vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__xor2_2
Xhold719 hold719/A vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14287_ _15448_/CLK hold980/X vssd1 vssd1 vccd1 vccd1 hold979/A sky130_fd_sc_hd__dfxtp_1
X_11499_ _11493_/A _11498_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _11499_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ _15357_/Q _15356_/Q _15355_/Q _15354_/Q vssd1 vssd1 vccd1 vccd1 _13239_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10173__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11984__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _13171_/A _13169_/B vssd1 vssd1 vccd1 vccd1 _15034_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2109 _14465_/Q vssd1 vssd1 vccd1 vccd1 hold2109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1408 _11911_/X vssd1 vssd1 vccd1 vccd1 _14732_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _14257_/Q vssd1 vssd1 vccd1 vccd1 hold1419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07730_ hold1553/X _13736_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07730_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__A2 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ hold1821/X _13700_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 _07661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_205_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09400_ _09400_/A _09400_/B vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12058__A0 hold2542/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13704__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07592_ _13698_/A1 hold2069/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07702__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ _09328_/Y _09329_/X _09161_/Y _09164_/Y vssd1 vssd1 vccd1 vccd1 _09331_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _09846_/B _10002_/C _09724_/C _09724_/D vssd1 vssd1 vccd1 vccd1 _09449_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__10084__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08213_ _09008_/A _08926_/A _08297_/A _08212_/D vssd1 vssd1 vccd1 vccd1 _08214_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ _09324_/A _09191_/Y _09060_/A _09060_/Y vssd1 vssd1 vccd1 vccd1 _09194_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09226__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08144_ _08144_/A _08144_/B _08144_/C vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_133_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07938__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12781__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _08892_/A _08075_/B _10507_/A _11550_/A vssd1 vssd1 vccd1 vccd1 _08077_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1076_A _13481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07026_ hold2021/X _13664_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07026_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08737__B1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11894__S _11894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06988__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2610 _15003_/Q vssd1 vssd1 vccd1 vccd1 hold2610/X sky130_fd_sc_hd__clkbuf_2
Xhold2621 _14978_/Q vssd1 vssd1 vccd1 vccd1 hold2621/X sky130_fd_sc_hd__buf_2
XANTENNA__13394__B _13394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2632 _15460_/Q vssd1 vssd1 vccd1 vccd1 hold2632/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _08989_/A _08976_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08977_/X sky130_fd_sc_hd__o21a_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout762_A _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2643 _09785_/X vssd1 vssd1 vccd1 vccd1 _14444_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2654 _12145_/X vssd1 vssd1 vccd1 vccd1 _14883_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2665 _14814_/Q vssd1 vssd1 vccd1 vccd1 hold2665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1920 _07154_/X vssd1 vssd1 vccd1 vccd1 _13962_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2676 _14813_/Q vssd1 vssd1 vccd1 vccd1 hold2676/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ hold203/A hold403/A hold971/A _13961_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07928_/X sky130_fd_sc_hd__mux4_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1931 _13987_/Q vssd1 vssd1 vccd1 vccd1 hold1931/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1942 _07100_/X vssd1 vssd1 vccd1 vccd1 _13913_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2687 _15139_/Q vssd1 vssd1 vccd1 vccd1 hold2687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2698 _14836_/Q vssd1 vssd1 vccd1 vccd1 hold2698/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1953 _13826_/Q vssd1 vssd1 vccd1 vccd1 hold1953/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1964 _07767_/X vssd1 vssd1 vccd1 vccd1 _14383_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1975 _14386_/Q vssd1 vssd1 vccd1 vccd1 hold1975/X sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _07859_/A vssd1 vssd1 vccd1 vccd1 _07859_/Y sky130_fd_sc_hd__inv_2
Xhold1986 _07753_/X vssd1 vssd1 vccd1 vccd1 _14369_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08060__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1997 _13868_/Q vssd1 vssd1 vccd1 vccd1 hold1997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10942__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _10870_/A _10870_/B vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07612__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09529_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09530_/C sky130_fd_sc_hd__a21bo_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ hold925/X hold1453/X _12665_/S vssd1 vssd1 vccd1 vccd1 _12540_/X sky130_fd_sc_hd__mux2_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12471_ _15364_/Q _15267_/Q _15075_/Q _14368_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12471_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_191_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12447__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _15398_/CLK hold496/X vssd1 vssd1 vccd1 vccd1 hold495/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ _11177_/B _11179_/B _11420_/X _11421_/Y vssd1 vssd1 vccd1 vccd1 _11449_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_117_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15190_ _15190_/CLK _15190_/D vssd1 vssd1 vccd1 vccd1 _15190_/Q sky130_fd_sc_hd__dfxtp_2
X_14141_ _15361_/CLK hold360/X vssd1 vssd1 vccd1 vccd1 hold359/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11353_ _11517_/A _15222_/Q _11352_/C _11352_/D vssd1 vssd1 vccd1 vccd1 _11354_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10783__B1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07059__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _11605_/A _11168_/A _10304_/C _10304_/D vssd1 vssd1 vccd1 vccd1 _10306_/D
+ sky130_fd_sc_hd__nand4_1
X_14072_ _15351_/CLK _14072_/D vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__dfxtp_1
X_11284_ _10955_/A _10955_/B _07318_/A vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ hold259/X hold317/A hold703/X _13986_/Q _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _13023_/X sky130_fd_sc_hd__mux4_1
X_10235_ _13750_/A _13365_/B _10233_/X _10234_/Y vssd1 vssd1 vccd1 vccd1 _10235_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12219__A_N _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ _10166_/A _10338_/B _10166_/C _10338_/C vssd1 vssd1 vccd1 vccd1 _10343_/A
+ sky130_fd_sc_hd__and4_1
X_14974_ _15004_/CLK hold160/X vssd1 vssd1 vccd1 vccd1 _14974_/Q sky130_fd_sc_hd__dfxtp_1
X_10097_ _14289_/Q _14225_/Q hold645/A _14479_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _10098_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12383__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13925_ _15458_/CLK _13925_/D vssd1 vssd1 vccd1 vccd1 _13925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08051__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13524__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ _14791_/CLK _13856_/D vssd1 vssd1 vccd1 vccd1 _13856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07522__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _13107_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _14960_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13787_ hold227/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__clkbuf_1
X_10999_ _10996_/Y _10997_/X _10793_/X _10816_/X vssd1 vssd1 vccd1 vccd1 _11033_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12917_/B1 _12733_/X _12737_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12745_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11979__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09208__A1 _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15457_ _15457_/CLK hold400/X vssd1 vssd1 vccd1 vccd1 hold399/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12669_ _12669_/A1 _12664_/X _12668_/X _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12670_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13004__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14408_ _15191_/CLK _14408_/D vssd1 vssd1 vccd1 vccd1 _14408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388_ _15457_/CLK hold954/X vssd1 vssd1 vccd1 vccd1 hold953/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09676__C _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12763__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14339_ _15436_/CLK hold500/X vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__dfxtp_1
Xhold505 hold505/A vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 hold516/A vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold527 hold527/A vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 hold538/A vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09973__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 hold549/A vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _08900_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _08901_/C sky130_fd_sc_hd__xor2_1
XANTENNA_hold2525_A _15353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _09879_/B _10030_/B _09879_/A vssd1 vssd1 vccd1 vccd1 _09881_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08721_/B _08721_/Y _08829_/Y _08830_/X vssd1 vssd1 vccd1 vccd1 _08948_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _14507_/Q vssd1 vssd1 vccd1 vccd1 hold1205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _11868_/X vssd1 vssd1 vccd1 vccd1 _14690_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08981_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _08762_/Y sky130_fd_sc_hd__nor2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 _14633_/Q vssd1 vssd1 vccd1 vccd1 hold1227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _06998_/X vssd1 vssd1 vccd1 vccd1 _13817_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1249 _14664_/Q vssd1 vssd1 vccd1 vccd1 hold1249/X sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ hold525/X _13719_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold526/A sky130_fd_sc_hd__mux2_1
X_08693_ _08694_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _08693_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07644_ _07644_/A _13683_/A vssd1 vssd1 vccd1 vccd1 _07644_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_164_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09790__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ _13404_/A _07575_/B vssd1 vssd1 vccd1 vccd1 _14200_/D sky130_fd_sc_hd__and2_1
XFILLER_0_211_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09314_ _09314_/A _09314_/B _09314_/C vssd1 vssd1 vccd1 vccd1 _09314_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08655__C1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11889__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _13734_/A1 _11514_/A2 _11514_/B1 _13189_/B _09243_/Y vssd1 vssd1 vccd1 vccd1
+ _09245_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout510_A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout608_A _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09176_ _09175_/B _09175_/C _09175_/A vssd1 vssd1 vccd1 vccd1 _09178_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13389__B _13389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12754__A1 _09342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08127_ _08201_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _08127_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10094__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08058_ _08065_/A _08055_/X _08057_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08059_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12506__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _13681_/A1 hold1019/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07009_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10822__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10020_ _10020_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07607__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput103 in1[15] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__clkbuf_1
Xinput114 in1[25] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_1
Xinput125 in1[6] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08281__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput136 in2[16] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__clkbuf_2
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2440 _12167_/X vssd1 vssd1 vccd1 vccd1 _14894_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2451 _15113_/Q vssd1 vssd1 vccd1 vccd1 hold2451/X sky130_fd_sc_hd__buf_1
Xinput147 in2[26] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__clkbuf_2
Xinput158 in2[7] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__clkbuf_2
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2462 _12117_/X vssd1 vssd1 vccd1 vccd1 _14870_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13467__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2473 _14450_/Q vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__buf_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2484 _12127_/X vssd1 vssd1 vccd1 vccd1 _14875_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2495 _14850_/Q vssd1 vssd1 vccd1 vccd1 hold2495/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12365__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1750 _07158_/X vssd1 vssd1 vccd1 vccd1 _13966_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1761 _13820_/Q vssd1 vssd1 vccd1 vccd1 hold1761/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ hold665/X _13512_/A0 _11977_/S vssd1 vssd1 vccd1 vccd1 hold666/A sky130_fd_sc_hd__mux2_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1772 _11714_/X vssd1 vssd1 vccd1 vccd1 _14510_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1783 _14377_/Q vssd1 vssd1 vccd1 vccd1 hold1783/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1794 _07098_/X vssd1 vssd1 vccd1 vccd1 _13911_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13710_ hold819/X _13743_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold820/A sky130_fd_sc_hd__mux2_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ _11108_/B _10749_/B _10745_/B vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__o21a_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _14754_/CLK _14690_/D vssd1 vssd1 vccd1 vccd1 _14690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _08253_/A _13625_/C _13640_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15353_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10853_ _10850_/X _10851_/Y _10631_/B _10633_/B vssd1 vssd1 vccd1 vccd1 _10853_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_116_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08646__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _14442_/Q _13590_/B vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__or2_1
XFILLER_0_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10784_ _11577_/A _11596_/A _14966_/Q vssd1 vssd1 vccd1 vccd1 _10784_/X sky130_fd_sc_hd__and3_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11799__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15311_ _15313_/CLK _15311_/D vssd1 vssd1 vccd1 vccd1 _15311_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12993__A1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ hold219/A _14306_/Q _14597_/Q _13966_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12523_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15242_ _15242_/CLK hold108/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_12454_ _13379_/B _12325_/B _12453_/X vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ _11158_/A _11158_/C _11158_/B vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07297__B _14964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15173_ _15177_/CLK _15173_/D vssd1 vssd1 vccd1 vccd1 _15173_/Q sky130_fd_sc_hd__dfxtp_2
X_12385_ hold957/A _13929_/Q _12460_/S vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__mux2_1
X_14124_ _15374_/CLK _14124_/D vssd1 vssd1 vccd1 vccd1 _14124_/Q sky130_fd_sc_hd__dfxtp_1
X_11336_ _11336_/A _11336_/B vssd1 vssd1 vccd1 vccd1 _11339_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13519__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _15340_/CLK _14055_/D vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__dfxtp_1
X_11267_ _11267_/A1 _11265_/X _11082_/A _11086_/A vssd1 vssd1 vccd1 vccd1 _11269_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10508__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09374__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ _13081_/A1 _13167_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _13007_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_197_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10218_ _10263_/C _10267_/A vssd1 vssd1 vccd1 vccd1 _10220_/C sky130_fd_sc_hd__nor2_1
X_11198_ _11195_/X _11382_/B _11006_/X _11009_/X vssd1 vssd1 vccd1 vccd1 _11199_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__A1 _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10149_ _10148_/B _10148_/C _10148_/A vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09677__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14957_ _14971_/CLK _14957_/D vssd1 vssd1 vccd1 vccd1 _14957_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11563__A _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ _15441_/CLK _13908_/D vssd1 vssd1 vccd1 vccd1 _13908_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12681__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14888_ _14889_/CLK _14888_/D vssd1 vssd1 vccd1 vccd1 _14888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09429__A1 _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__A _14941_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13839_ _15391_/CLK _13839_/D vssd1 vssd1 vccd1 vccd1 _13839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09429__B2 _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07360_ _07362_/B _07360_/B _07353_/C vssd1 vssd1 vccd1 vccd1 _07360_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07291_ _11542_/B _10115_/D vssd1 vssd1 vccd1 vccd1 _09767_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09030_ _09030_/A _09030_/B _09030_/C vssd1 vssd1 vccd1 vccd1 _09032_/A sky130_fd_sc_hd__and3_1
XFILLER_0_14_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__A2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10747__B1 _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold313 hold313/A vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 hold346/A vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold357 hold357/A vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09932_ _10401_/A _09932_/B _09932_/C vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__and3_1
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 hold379/A vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10642__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout804 _12365_/S1 vssd1 vssd1 vccd1 vccd1 _12689_/S1 sky130_fd_sc_hd__buf_8
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout815 _14489_/Q vssd1 vssd1 vccd1 vccd1 _13068_/A1 sky130_fd_sc_hd__buf_2
Xfanout826 _12560_/S vssd1 vssd1 vccd1 vccd1 _12665_/S sky130_fd_sc_hd__buf_6
X_09863_ _09864_/A _10022_/A _10304_/C _10304_/D vssd1 vssd1 vccd1 vccd1 _09863_/X
+ sky130_fd_sc_hd__and4_1
Xfanout837 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _13066_/S sky130_fd_sc_hd__buf_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout848 _13481_/A vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__clkbuf_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout859 _07473_/B vssd1 vssd1 vccd1 vccd1 _13622_/C1 sky130_fd_sc_hd__clkbuf_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08814_/A _08814_/B _08814_/C vssd1 vssd1 vccd1 vccd1 _08816_/B sky130_fd_sc_hd__nand3_2
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _07008_/X vssd1 vssd1 vccd1 vccd1 _13827_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _15368_/Q vssd1 vssd1 vccd1 vccd1 hold1013/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _10246_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _09794_/Y sky130_fd_sc_hd__nor2_1
Xhold1024 _13657_/X vssd1 vssd1 vccd1 vccd1 _15364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 _13814_/Q vssd1 vssd1 vccd1 vccd1 hold1035/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1046 _07068_/X vssd1 vssd1 vccd1 vccd1 _13884_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08642_/A _08642_/B _08639_/X vssd1 vssd1 vccd1 vccd1 _08746_/B sky130_fd_sc_hd__a21o_1
Xhold1057 _14631_/Q vssd1 vssd1 vccd1 vccd1 hold1057/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 _11749_/X vssd1 vssd1 vccd1 vccd1 _14543_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1079 _14422_/Q vssd1 vssd1 vccd1 vccd1 hold1079/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12898__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11473__A _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__A1 _07879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_208 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08676_ _08901_/A _08892_/A _09866_/B _09864_/C vssd1 vssd1 vccd1 vccd1 _08785_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA_219 _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07162__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12288__B _12288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07627_ hold545/X _13700_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold546/A sky130_fd_sc_hd__mux2_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout725_A _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09878__A _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _13393_/A hold149/X vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__and2_1
XANTENNA__09515__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14934__D _14934_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07489_ hold1851/X _13728_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07489_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ hold373/A _15278_/Q hold347/A _14379_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09228_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13075__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ _09159_/A _09159_/B vssd1 vssd1 vccd1 vccd1 _09160_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10738__B1 _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07829__S1 _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12170_ _14896_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11121_ _11497_/A _11120_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _11121_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold880 hold880/A vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 hold891/A vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__xor2_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10271__B _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10005_/B sky130_fd_sc_hd__nor2_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2270 _11926_/X vssd1 vssd1 vccd1 vccd1 _14747_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07861__A _15345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12338__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2281 _15329_/Q vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13582__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ _15196_/CLK _14811_/D vssd1 vssd1 vccd1 vccd1 _14811_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2292 _07156_/X vssd1 vssd1 vccd1 vccd1 _13964_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08676__B _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12889__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1580 _11773_/X vssd1 vssd1 vccd1 vccd1 _14598_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11954_ _13742_/A1 hold2159/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11954_/X sky130_fd_sc_hd__mux2_1
X_14742_ _15242_/CLK _14742_/D vssd1 vssd1 vccd1 vccd1 _14742_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1591 _13895_/Q vssd1 vssd1 vccd1 vccd1 hold1591/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07072__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _11091_/A _10903_/Y _10717_/B _10719_/C vssd1 vssd1 vccd1 vccd1 _10905_/X
+ sky130_fd_sc_hd__o211a_1
X_14673_ _15448_/CLK _14673_/D vssd1 vssd1 vccd1 vccd1 _14673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ hold491/X _13739_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold492/A sky130_fd_sc_hd__mux2_1
XANTENNA__15005__D _15005_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13624_ _08849_/A _13792_/A2 _13623_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15339_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ _10836_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07800__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ _08435_/B _08441_/B _13554_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _15303_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10767_ _11493_/A _10767_/B vssd1 vssd1 vccd1 vccd1 _10767_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_171_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08634__A2 _13385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _08253_/A _08636_/A _13147_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12507_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12420__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__B _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13486_ _13486_/A hold121/X vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__and2_1
X_10698_ _14947_/Q _11561_/A _11542_/B _11564_/B vssd1 vssd1 vccd1 vccd1 _10878_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_125_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12718__A1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15225_ _15225_/CLK _15225_/D vssd1 vssd1 vccd1 vccd1 _15225_/Q sky130_fd_sc_hd__dfxtp_2
X_12437_ _12674_/S1 _12434_/X _12436_/X vssd1 vssd1 vccd1 vccd1 _12437_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _15423_/CLK _15156_/D vssd1 vssd1 vccd1 vccd1 _15156_/Q sky130_fd_sc_hd__dfxtp_1
X_12368_ _12368_/A _12368_/B vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__and2_1
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12570__C_N _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ _15360_/CLK hold896/X vssd1 vssd1 vccd1 vccd1 hold895/A sky130_fd_sc_hd__dfxtp_1
X_11319_ _11304_/Y _11309_/Y _11318_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _11320_/B sky130_fd_sc_hd__a221o_1
X_15087_ _15087_/CLK hold690/X vssd1 vssd1 vccd1 vccd1 hold689/A sky130_fd_sc_hd__dfxtp_1
X_12299_ _15346_/Q _07875_/C _07875_/B _15347_/Q vssd1 vssd1 vccd1 vccd1 _12299_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14038_ _14083_/CLK _14038_/D vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12351__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08530_ _08530_/A _08530_/B _08530_/C _08530_/D vssd1 vssd1 vccd1 vccd1 _08530_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08461_ hold199/A _14535_/Q hold429/A _14759_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08461_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_187_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_183_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _14397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07412_ _13501_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _14042_/D sky130_fd_sc_hd__and2_1
XANTENNA__13712__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__B1 _13143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08393_/A _08393_/B _08393_/C vssd1 vssd1 vccd1 vccd1 _08392_/X sky130_fd_sc_hd__and3_1
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07343_ _14059_/Q _14060_/Q _14062_/Q _14063_/Q vssd1 vssd1 vccd1 vccd1 _07343_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_175_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10637__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07274_ _07274_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08107__A _08107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _08892_/X _08894_/X _09011_/Y _09012_/X vssd1 vssd1 vccd1 vccd1 _09013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12852__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _09860_/B vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07157__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _15207_/Q vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__clkbuf_8
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _09914_/A _09914_/C _09914_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__a21o_1
Xfanout623 _15204_/Q vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__clkbuf_8
Xfanout634 _15201_/Q vssd1 vssd1 vccd1 vccd1 _11597_/A sky130_fd_sc_hd__clkbuf_8
Xfanout645 _15199_/Q vssd1 vssd1 vccd1 vccd1 _10002_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout675_A _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout656 _13681_/A1 vssd1 vssd1 vccd1 vccd1 _13714_/A1 sky130_fd_sc_hd__clkbuf_4
X_09846_ _10000_/A _09846_/B _11605_/B _10108_/C vssd1 vssd1 vccd1 vccd1 _10005_/A
+ sky130_fd_sc_hd__and4_1
Xfanout667 _15062_/Q vssd1 vssd1 vccd1 vccd1 _13742_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06996__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout678 _13704_/A1 vssd1 vssd1 vccd1 vccd1 _13737_/A1 sky130_fd_sc_hd__buf_2
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _15052_/Q vssd1 vssd1 vccd1 vccd1 _13732_/A1 sky130_fd_sc_hd__buf_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14929__D _14929_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _09218_/A _09349_/A _09491_/A _09628_/A _09776_/X vssd1 vssd1 vccd1 vccd1
+ _09930_/A sky130_fd_sc_hd__o41a_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _13661_/A1 hold1537/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06989_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout842_A _14488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08728_ _08725_/X _08726_/Y _08593_/X _08596_/X vssd1 vssd1 vccd1 vccd1 _08728_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08313__A1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ hold611/A _14214_/Q hold555/A _14468_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08660_/B sky130_fd_sc_hd__mux4_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15177_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11670_ _13734_/A1 hold873/X _11684_/S vssd1 vssd1 vccd1 vccd1 hold874/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10621_ _11597_/A _11598_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _10623_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _13342_/A _13340_/B vssd1 vssd1 vccd1 vccd1 _13750_/B sky130_fd_sc_hd__or2_1
X_10552_ _10553_/A _10553_/B _10553_/C vssd1 vssd1 vccd1 vccd1 _10552_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13048__S1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ input96/X fanout1/X _13270_/X vssd1 vssd1 vccd1 vccd1 _13272_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ _10483_/A _10483_/B vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15010_ _15177_/CLK _15010_/D vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__dfxtp_1
X_12222_ _12221_/B _12220_/X _12221_/Y vssd1 vssd1 vccd1 vccd1 _13374_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09041__A2 _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ hold2617/X _12173_/A2 _12152_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07067__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ _11104_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _11104_/X sky130_fd_sc_hd__and2_1
XFILLER_0_208_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12084_ _14982_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12084_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_159_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11035_ _11035_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11037_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__B1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ _13092_/A1 _12985_/X _13050_/S0 vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08304__A1 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__B2 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14725_ _14783_/CLK _14725_/D vssd1 vssd1 vccd1 vccd1 _14725_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__A1 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ _13725_/A1 hold1137/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_165_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15405_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13532__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14656_ _15434_/CLK hold958/X vssd1 vssd1 vccd1 vccd1 hold957/A sky130_fd_sc_hd__dfxtp_1
X_11868_ hold1215/X _13689_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07530__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _10819_/A _10819_/B _10819_/C vssd1 vssd1 vccd1 vccd1 _11037_/A sky130_fd_sc_hd__nand3_2
X_13607_ input60/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13607_/X sky130_fd_sc_hd__or2_1
XFILLER_0_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13061__B1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14587_ _14651_/CLK hold214/X vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__dfxtp_1
X_11799_ hold763/X _13653_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold764/A sky130_fd_sc_hd__mux2_1
XANTENNA__13600__A2 _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13538_ _15460_/Q _13634_/B vssd1 vssd1 vccd1 vccd1 _13538_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13039__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11987__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13469_ _11645_/B _13468_/A _13468_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 _13469_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15226_/CLK _15208_/D vssd1 vssd1 vccd1 vccd1 _15208_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12798__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput204 _14187_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[17] sky130_fd_sc_hd__buf_12
XFILLER_0_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput215 _14197_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[27] sky130_fd_sc_hd__buf_12
XFILLER_0_140_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput226 _14178_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[8] sky130_fd_sc_hd__buf_12
Xoutput237 _14442_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[18] sky130_fd_sc_hd__buf_12
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput248 _14452_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[28] sky130_fd_sc_hd__buf_12
XFILLER_0_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15139_ _15299_/CLK _15139_/D vssd1 vssd1 vccd1 vccd1 _15139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput259 _14433_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[9] sky130_fd_sc_hd__buf_12
XFILLER_0_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09981__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _07961_/A _07961_/B vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11438__D _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _09702_/D vssd1 vssd1 vccd1 vccd1 _09700_/Y sky130_fd_sc_hd__inv_2
X_06912_ _15341_/Q vssd1 vssd1 vccd1 vccd1 _07862_/C sky130_fd_sc_hd__inv_2
XANTENNA__13707__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2605_A _14994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07892_ _08677_/A _10873_/A _08892_/A _08312_/A vssd1 vssd1 vccd1 vccd1 _07894_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__10920__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07705__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _09499_/X _09630_/X _13586_/B vssd1 vssd1 vccd1 vccd1 _09631_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13419__A2 _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09562_ _09846_/B _10283_/C _10115_/D _10000_/A vssd1 vssd1 vccd1 vccd1 _09562_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08513_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_195_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12722__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10102__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _09918_/A _13442_/B _13360_/B _08256_/A _09492_/Y vssd1 vssd1 vccd1 vccd1
+ _09493_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_210_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_156_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15391_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ _08542_/A _08544_/C vssd1 vssd1 vccd1 vccd1 _08444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10653__A2 _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ hold2745/X input32/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13181_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout423_A _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07326_ _07326_/A _10956_/A _07326_/C _07326_/D vssd1 vssd1 vccd1 vccd1 _07329_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_128_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11897__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07257_ _11168_/A _10304_/C vssd1 vssd1 vccd1 vccd1 _07258_/B sky130_fd_sc_hd__or2_1
XFILLER_0_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12789__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13397__B _13397_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07188_ hold387/X _13656_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold388/A sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08457__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout420 _13650_/Y vssd1 vssd1 vccd1 vccd1 _13682_/S sky130_fd_sc_hd__buf_12
Xfanout431 _11763_/Y vssd1 vssd1 vccd1 vccd1 _11779_/S sky130_fd_sc_hd__buf_12
XFILLER_0_10_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07990__C1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 _07389_/Y vssd1 vssd1 vccd1 vccd1 _08441_/B sky130_fd_sc_hd__buf_4
Xfanout453 _13636_/B vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__buf_2
Xfanout464 _07045_/X vssd1 vssd1 vccd1 vccd1 _07077_/S sky130_fd_sc_hd__clkbuf_16
Xfanout475 _13466_/A vssd1 vssd1 vccd1 vccd1 _13468_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07615__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09829_ _09709_/D _09711_/A _09827_/Y _09828_/X vssd1 vssd1 vccd1 vccd1 _09831_/B
+ sky130_fd_sc_hd__a211o_2
Xfanout497 _06943_/Y vssd1 vssd1 vccd1 vccd1 _12669_/A1 sky130_fd_sc_hd__buf_8
X_12840_ hold1127/X _14127_/Q _12841_/S vssd1 vssd1 vccd1 vccd1 _12840_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_198_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12771_ _15376_/Q _15279_/Q hold689/A _14380_/Q _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12771_/X sky130_fd_sc_hd__mux4_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_147_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _14775_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14510_ _15188_/CLK _14510_/D vssd1 vssd1 vccd1 vccd1 _14510_/Q sky130_fd_sc_hd__dfxtp_1
X_11722_ hold431/X _11921_/A0 _11728_/S vssd1 vssd1 vccd1 vccd1 hold432/A sky130_fd_sc_hd__mux2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__A2 _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__B _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _15313_/CLK _14441_/D vssd1 vssd1 vccd1 vccd1 _14441_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _12329_/A hold1201/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ _11580_/A _14967_/Q vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__nand2_1
X_14372_ _15079_/CLK _14372_/D vssd1 vssd1 vccd1 vccd1 _14372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13323_ _13338_/A _13323_/B vssd1 vssd1 vccd1 vccd1 _15127_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_181_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10535_ _10534_/B _10534_/C _10534_/A vssd1 vssd1 vccd1 vccd1 _10535_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_107_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08470__B1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ _13287_/A _13254_/B vssd1 vssd1 vccd1 vccd1 _15104_/D sky130_fd_sc_hd__nor2_1
X_10466_ _10635_/A _10467_/C _10467_/A vssd1 vssd1 vccd1 vccd1 _10502_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output175_A _15186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _12233_/A _12204_/X _12247_/A vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13185_ _13393_/A _13185_/B vssd1 vssd1 vccd1 vccd1 _15050_/D sky130_fd_sc_hd__and2_1
X_10397_ _10397_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10397_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_209_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _14879_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12136_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10580__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13527__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12067_ hold2487/X _12099_/A2 _12066_/X _13492_/A vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09948__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07525__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11018_ _09075_/A _11018_/B _11201_/A vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08210__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15449_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _13100_/S0 _12964_/X _12968_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _12970_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14708_ _15450_/CLK hold326/X vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _15087_/CLK _14639_/D vssd1 vssd1 vccd1 vccd1 _14639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13585__A1 _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08160_ _08289_/A _08159_/B _08093_/A vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_32_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ _13714_/A1 hold2181/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13498__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _08091_/A _08091_/B vssd1 vssd1 vccd1 vccd1 _08093_/C sky130_fd_sc_hd__and2_1
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2555_A _14998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07042_ hold945/X _13680_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold946/A sky130_fd_sc_hd__mux2_1
XFILLER_0_140_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07016__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _08978_/Y _08983_/Y _08992_/X _12241_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08994_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2803 _13895_/Q vssd1 vssd1 vccd1 vccd1 hold2803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2814 _14114_/Q vssd1 vssd1 vccd1 vccd1 hold2814/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold2825 _15325_/Q vssd1 vssd1 vccd1 vccd1 hold2825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07944_ _08197_/A _07943_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _07944_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2836 _15339_/Q vssd1 vssd1 vccd1 vccd1 hold2836/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09939__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2847 _15308_/Q vssd1 vssd1 vccd1 vccd1 hold2847/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2858 _14022_/Q vssd1 vssd1 vccd1 vccd1 hold2858/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07875_ _11763_/B _07875_/B _07875_/C vssd1 vssd1 vccd1 vccd1 _07875_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_39_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09614_ _09760_/B _09759_/D vssd1 vssd1 vccd1 vccd1 _09616_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09545_ _09545_/A _09673_/B _09545_/C vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_leaf_129_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15377_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout540_A _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12577__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _15200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ _09202_/A _09335_/A _09333_/X vssd1 vssd1 vccd1 vccd1 _09476_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07170__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08427_ _08519_/B _08427_/B _08427_/C vssd1 vssd1 vccd1 vccd1 _08428_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_114_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_A _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08358_ _08873_/A _08355_/X _08357_/X vssd1 vssd1 vccd1 vccd1 _08358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_191_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08790__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07309_ _07324_/A vssd1 vssd1 vccd1 vccd1 _08172_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08289_ _08289_/A _08326_/B vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__and2_1
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12516__S _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13328__A1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ _10320_/A _10320_/B _10320_/C vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13201__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ hold771/A _13950_/Q hold355/A _13918_/Q _10425_/S0 _10425_/S1 vssd1 vssd1
+ vccd1 vccd1 _10252_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08755__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10182_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10189_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_206_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14990_ _15248_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 _14990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11375__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13941_ _15439_/CLK _13941_/D vssd1 vssd1 vccd1 vccd1 _13941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08387__D _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13872_ _15079_/CLK _13872_/D vssd1 vssd1 vccd1 vccd1 _13872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12823_ hold207/A _14318_/Q _14609_/Q _13978_/Q _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12823_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13590__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08366__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12754_ _09342_/X _13104_/A2 _12753_/X vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__a21o_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ hold709/X _13659_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold710/A sky130_fd_sc_hd__mux2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _14668_/Q _13941_/Q _12735_/S vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15013__D _15013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11636_ _11636_/A _11636_/B vssd1 vssd1 vccd1 vccd1 _11637_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09796__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14424_ _15068_/CLK hold474/X vssd1 vssd1 vccd1 vccd1 hold473/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11567_/A _15228_/Q vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__nand2_1
X_14355_ _15383_/CLK _14355_/D vssd1 vssd1 vccd1 vccd1 _14355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09640__C1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13319__A1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ input142/X fanout5/X fanout3/X input110/X vssd1 vssd1 vccd1 vccd1 _13306_/X
+ sky130_fd_sc_hd__a22o_1
X_10518_ _11340_/A _15220_/Q _10347_/A _10344_/X vssd1 vssd1 vccd1 vccd1 _10519_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14286_ _15410_/CLK hold806/X vssd1 vssd1 vccd1 vccd1 hold805/A sky130_fd_sc_hd__dfxtp_1
Xhold709 hold709/A vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11498_ _15421_/Q _14556_/Q hold571/A _14780_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11498_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13237_ _15351_/Q _15350_/Q vssd1 vssd1 vccd1 vccd1 _13239_/C sky130_fd_sc_hd__nor2_1
X_10449_ _11597_/A _11569_/B _11563_/B _11596_/A vssd1 vssd1 vccd1 vccd1 _10450_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_161_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _13168_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _15033_/D sky130_fd_sc_hd__nor2_1
XANTENNA__09962__C _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12119_ hold2493/X _12129_/A2 _12118_/X _13501_/A vssd1 vssd1 vccd1 vccd1 _12119_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_41_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ _13893_/Q _14021_/Q hold871/A _13829_/Q _13091_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13099_/X sky130_fd_sc_hd__mux4_1
Xhold1409 _13829_/Q vssd1 vssd1 vccd1 vccd1 hold1409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09036__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12925__S0 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_176_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ hold757/X _13732_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold758/A sky130_fd_sc_hd__mux2_1
XANTENNA__08875__A _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_56_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07591_ _13730_/A1 hold1143/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07591_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09330_ _09161_/Y _09164_/Y _09328_/Y _09329_/X vssd1 vssd1 vccd1 vccd1 _09330_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10001__A1_N _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09261_ _10002_/C _09724_/C _09724_/D _09846_/B vssd1 vssd1 vccd1 vccd1 _09264_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08212_ _09008_/A _08926_/A _08297_/A _08212_/D vssd1 vssd1 vccd1 vccd1 _08297_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__13720__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ _09060_/A _09060_/Y _09324_/A _09191_/Y vssd1 vssd1 vccd1 vccd1 _09328_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08143_ _08776_/A _10507_/A _11550_/A _09008_/A vssd1 vssd1 vccd1 vccd1 _08144_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10645__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08074_ _11566_/A _08776_/A vssd1 vssd1 vccd1 vccd1 _08077_/A sky130_fd_sc_hd__and2_1
XANTENNA__12781__A2 _13158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07025_ hold1879/X _13663_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07025_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_129_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11476__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2600 hold2861/X vssd1 vssd1 vccd1 vccd1 hold2600/X sky130_fd_sc_hd__buf_1
Xhold2611 _12193_/X vssd1 vssd1 vccd1 vccd1 _14907_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2622 _12143_/X vssd1 vssd1 vccd1 vccd1 _14882_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08976_ _13877_/Q hold713/A _13845_/Q _13813_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08976_/X sky130_fd_sc_hd__mux4_1
Xhold2633 _13755_/X vssd1 vssd1 vccd1 vccd1 _15460_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2644 _14437_/Q vssd1 vssd1 vccd1 vccd1 _08856_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1910 _11784_/X vssd1 vssd1 vccd1 vccd1 _14609_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2655 _15330_/Q vssd1 vssd1 vccd1 vccd1 hold2655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2666 _12002_/X vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1921 _14137_/Q vssd1 vssd1 vccd1 vccd1 hold1921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _07924_/X _07926_/Y _13369_/A vssd1 vssd1 vccd1 vccd1 _07927_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2677 _12000_/X vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1932 _07179_/X vssd1 vssd1 vccd1 vccd1 _13987_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A _14950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2688 _08184_/Y vssd1 vssd1 vccd1 vccd1 hold2688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1943 _13959_/Q vssd1 vssd1 vccd1 vccd1 hold1943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2699 _14840_/Q vssd1 vssd1 vccd1 vccd1 hold2699/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1954 _07007_/X vssd1 vssd1 vccd1 vccd1 _13826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1965 _13949_/Q vssd1 vssd1 vccd1 vccd1 hold1965/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07858_ _07341_/B _07847_/X _07857_/X _12256_/A _07885_/B vssd1 vssd1 vccd1 vccd1
+ _07859_/A sky130_fd_sc_hd__o311a_1
Xhold1976 _07770_/X vssd1 vssd1 vccd1 vccd1 _14386_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1987 _14385_/Q vssd1 vssd1 vccd1 vccd1 hold1987/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1998 _07052_/X vssd1 vssd1 vccd1 vccd1 _13868_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14937__D _14937_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07789_ hold959/X _13727_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold960/A sky130_fd_sc_hd__mux2_1
XFILLER_0_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09528_ _09527_/B _09527_/C _09527_/A vssd1 vssd1 vccd1 vccd1 _09530_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_151_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12100__A _14990_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08122__C1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _09459_/A _09599_/A _09459_/C vssd1 vssd1 vccd1 vccd1 _09461_/C sky130_fd_sc_hd__nand3_4
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _12470_/A _12470_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12477_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ _11551_/B _11420_/C _11420_/A vssd1 vssd1 vccd1 vccd1 _11421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14140_ _15392_/CLK _14140_/D vssd1 vssd1 vccd1 vccd1 _14140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _11517_/A _15222_/Q _11352_/C _11352_/D vssd1 vssd1 vccd1 vccd1 _11354_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08025__A _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10783__A1 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _11605_/A _11168_/A _11542_/A _11536_/A vssd1 vssd1 vccd1 vccd1 _10303_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10783__B2 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14071_ _15293_/CLK _14071_/D vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__dfxtp_1
X_11283_ hold2779/X _11282_/Y _11283_/S vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ hold371/X hold349/X hold363/X hold2009/X _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _13022_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09925__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _15156_/Q _07812_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _10234_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10165_ _10338_/B _10166_/C _10338_/C _10166_/A vssd1 vssd1 vccd1 vccd1 _10165_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__07075__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14973_ _14973_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 _14973_/Q sky130_fd_sc_hd__dfxtp_1
X_10096_ _11493_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10096_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12383__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _15457_/CLK _13924_/D vssd1 vssd1 vccd1 vccd1 _13924_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08695__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07803__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ _15415_/CLK hold740/X vssd1 vssd1 vccd1 vccd1 hold739/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12806_ _13106_/A1 _13159_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_174_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10998_ _10793_/X _10816_/X _10996_/Y _10997_/X vssd1 vssd1 vccd1 vccd1 _11033_/A
+ sky130_fd_sc_hd__o211ai_4
X_13786_ hold213/X vssd1 vssd1 vccd1 vccd1 hold214/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08113__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08664__B1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12749_/S1 _12734_/X _12736_/X vssd1 vssd1 vccd1 vccd1 _12737_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13540__S _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__C _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15456_ _15456_/CLK hold830/X vssd1 vssd1 vccd1 vccd1 hold829/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06943__A _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12668_ _12668_/A1 _12665_/X _12667_/X vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _14602_/CLK hold970/X vssd1 vssd1 vccd1 vccd1 hold969/A sky130_fd_sc_hd__dfxtp_1
X_11619_ _11454_/A _11453_/B _11453_/A vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15387_ _15387_/CLK _15387_/D vssd1 vssd1 vccd1 vccd1 _15387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09676__D _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ _13873_/Q hold891/A hold687/A _13809_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12599_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ _15437_/CLK hold462/X vssd1 vssd1 vccd1 vccd1 hold461/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold506 hold506/A vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10774__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 hold517/A vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold528 hold528/A vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09973__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold539 hold539/A vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14269_ _14397_/CLK hold424/X vssd1 vssd1 vccd1 vccd1 hold423/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08829_/B _08829_/C _08829_/A vssd1 vssd1 vccd1 vccd1 _08830_/X sky130_fd_sc_hd__o21a_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _11711_/X vssd1 vssd1 vccd1 vccd1 _14507_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 _14778_/Q vssd1 vssd1 vccd1 vccd1 hold1217/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ hold989/A _14247_/Q hold969/A _14119_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08762_/B sky130_fd_sc_hd__mux4_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _11809_/X vssd1 vssd1 vccd1 vccd1 _14633_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1239 _14135_/Q vssd1 vssd1 vccd1 vccd1 hold1239/X sky130_fd_sc_hd__dlygate4sd3_1
X_07712_ hold2155/X _13718_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 _07712_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13715__S _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11487__C1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ _08692_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07713__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07643_ _14086_/Q _14087_/Q _07643_/C _11763_/B vssd1 vssd1 vccd1 vccd1 _13683_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07574_ _13404_/A _07574_/B vssd1 vssd1 vccd1 vccd1 _14199_/D sky130_fd_sc_hd__and2_1
XFILLER_0_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _09314_/A _09314_/B _09314_/C vssd1 vssd1 vccd1 vccd1 _09317_/B sky130_fd_sc_hd__and3_1
XFILLER_0_165_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12581__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14842_/CLK sky130_fd_sc_hd__clkbuf_16
X_09244_ hold2738/X input9/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _09175_/A _09175_/B _09175_/C vssd1 vssd1 vccd1 vccd1 _09178_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout503_A _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08126_ _14272_/Q _14208_/Q _14144_/Q _14462_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08127_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12754__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08057_ _08981_/A _08057_/B vssd1 vssd1 vccd1 vccd1 _08057_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07008_ _13680_/A1 hold1001/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07008_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout872_A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput104 in1[16] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput115 in1[26] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11190__A1 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput126 in1[7] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_1
Xhold2430 _15312_/Q vssd1 vssd1 vccd1 vccd1 _06916_/A sky130_fd_sc_hd__buf_1
Xinput137 in2[17] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__clkbuf_2
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2441 _15131_/Q vssd1 vssd1 vccd1 vccd1 hold2441/X sky130_fd_sc_hd__buf_1
Xinput148 in2[27] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__clkbuf_2
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2452 _14849_/Q vssd1 vssd1 vccd1 vccd1 hold2452/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput159 in2[8] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__clkbuf_2
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ _07230_/A _08845_/X _07327_/B vssd1 vssd1 vccd1 vccd1 _09075_/C sky130_fd_sc_hd__a21o_1
Xhold2463 hold2846/X vssd1 vssd1 vccd1 vccd1 _08640_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2474 _10756_/X vssd1 vssd1 vccd1 vccd1 _14450_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1740 _07581_/X vssd1 vssd1 vccd1 vccd1 _14205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2485 _15000_/Q vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__buf_2
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1751 _13866_/Q vssd1 vssd1 vccd1 vccd1 hold1751/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12365__S1 _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2496 _12077_/X vssd1 vssd1 vccd1 vccd1 _14850_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1762 _07001_/X vssd1 vssd1 vccd1 vccd1 _13820_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11970_ hold1471/X _13659_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__mux2_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1773 _14680_/Q vssd1 vssd1 vccd1 vccd1 hold1773/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1784 _07761_/X vssd1 vssd1 vccd1 vccd1 _14377_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07623__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09404__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1795 _14756_/Q vssd1 vssd1 vccd1 vccd1 hold1795/X sky130_fd_sc_hd__dlygate4sd3_1
X_10921_ _11645_/A _10921_/B vssd1 vssd1 vccd1 vccd1 _11108_/D sky130_fd_sc_hd__xnor2_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13640_ input52/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13640_/X sky130_fd_sc_hd__or2_1
X_10852_ _10631_/B _10633_/B _10850_/X _10851_/Y vssd1 vssd1 vccd1 vccd1 _10852_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10783_ _11596_/A _11573_/B _14966_/Q _11577_/A vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12442__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _09346_/A _09222_/B _13570_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13571_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15340_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08110__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15310_ _15313_/CLK _15310_/D vssd1 vssd1 vccd1 vccd1 _15310_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _14789_/Q hold709/A hold375/A _14725_/Q _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12522_/X sky130_fd_sc_hd__mux4_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15241_ _15243_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12453_ _13656_/A1 _12329_/B _12953_/B1 _13177_/B vssd1 vssd1 vccd1 vccd1 _12453_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15172_ _15268_/CLK _15172_/D vssd1 vssd1 vccd1 vccd1 _15172_/Q sky130_fd_sc_hd__dfxtp_2
X_12384_ _15430_/Q _13897_/Q _12460_/S vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11953__A0 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11335_ _11335_/A _15225_/Q vssd1 vssd1 vccd1 vccd1 _11336_/B sky130_fd_sc_hd__nand2_1
X_14123_ _15375_/CLK _14123_/D vssd1 vssd1 vccd1 vccd1 _14123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11266_ _11082_/A _11086_/A _11267_/A1 _11265_/X vssd1 vssd1 vccd1 vccd1 _11465_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14054_ _15340_/CLK _14054_/D vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10508__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10508__B2 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output255_A _14429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ _10065_/B _10065_/Y _10392_/B _10215_/X vssd1 vssd1 vccd1 vccd1 _10267_/A
+ sky130_fd_sc_hd__a211oi_2
X_13005_ _13080_/A1 _13004_/X _13002_/X vssd1 vssd1 vccd1 vccd1 _13167_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11197_ _11006_/X _11009_/X _11195_/X _11382_/B vssd1 vssd1 vccd1 vccd1 _11197_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07924__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _10148_/A _10148_/B _10148_/C vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09126__A1 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10079_ _06940_/Y _12256_/A _10075_/X _10078_/X vssd1 vssd1 vccd1 vccd1 _13396_/B
+ sky130_fd_sc_hd__o211ai_4
X_14956_ _14956_/CLK _14956_/D vssd1 vssd1 vccd1 vccd1 _14956_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09677__A2 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11563__B _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _15440_/CLK _13907_/D vssd1 vssd1 vccd1 vccd1 _13907_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12681__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14887_ _14889_/CLK _14887_/D vssd1 vssd1 vccd1 vccd1 _14887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08980__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13838_ _14783_/CLK hold906/X vssd1 vssd1 vccd1 vccd1 hold905/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09429__A2 _14950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__B _15220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12969__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13769_ hold235/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _14105_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07290_ _09205_/B _07290_/B vssd1 vssd1 vccd1 vccd1 _09075_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_116_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15439_ _15439_/CLK hold956/X vssd1 vssd1 vccd1 vccd1 hold955/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11944__A0 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold314 hold314/A vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 hold336/A vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold347 hold347/A vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07708__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold358 hold358/A vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_09931_ _09932_/B _09932_/C _10401_/A vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__a21oi_1
Xhold369 hold369/A vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10642__B _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout805 _12365_/S1 vssd1 vssd1 vccd1 vccd1 _12343_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__09365__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout816 _13098_/S1 vssd1 vssd1 vccd1 vccd1 _13024_/S1 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_4_7__f_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09862_ _09712_/A _09864_/C _09864_/D _09864_/A vssd1 vssd1 vccd1 vccd1 _09866_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout827 _12560_/S vssd1 vssd1 vccd1 vccd1 _12566_/S sky130_fd_sc_hd__buf_6
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout838 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _12941_/S sky130_fd_sc_hd__buf_6
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _13477_/A vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__clkbuf_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _08922_/B _08812_/C _08812_/A vssd1 vssd1 vccd1 vccd1 _08814_/C sky130_fd_sc_hd__a21o_1
Xhold1003 _14139_/Q vssd1 vssd1 vccd1 vccd1 hold1003/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _10426_/A _09790_/X _09792_/X _10255_/A1 vssd1 vssd1 vccd1 vccd1 _09794_/B
+ sky130_fd_sc_hd__o211a_1
Xhold1014 _13661_/X vssd1 vssd1 vccd1 vccd1 _15368_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1025 _13835_/Q vssd1 vssd1 vccd1 vccd1 hold1025/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _06995_/X vssd1 vssd1 vccd1 vccd1 _13814_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 _15433_/Q vssd1 vssd1 vccd1 vccd1 hold1047/X sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _08742_/X _08744_/B vssd1 vssd1 vccd1 vccd1 _08746_/A sky130_fd_sc_hd__and2b_1
Xhold1058 _11807_/X vssd1 vssd1 vccd1 vccd1 _14631_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1069 _14469_/Q vssd1 vssd1 vccd1 vccd1 hold1069/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08893_/A _09866_/B _09864_/C _08677_/A vssd1 vssd1 vccd1 vccd1 _08678_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_209 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout453_A _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07626_ hold601/X _13732_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 hold602/A sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07557_ _13393_/A hold129/X vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__and2_1
XFILLER_0_49_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout620_A _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15435_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10435__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07488_ hold561/X _13727_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 hold562/A sky130_fd_sc_hd__mux2_1
XFILLER_0_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10986__A1 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09227_ _09941_/A _09224_/X _09226_/X vssd1 vssd1 vccd1 vccd1 _09227_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09158_ _09157_/A _09157_/B _09157_/C vssd1 vssd1 vccd1 vccd1 _09159_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08109_ _08109_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09089_ _10233_/A _09350_/C _09089_/C vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__or3_1
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07618__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120_ _13891_/Q _14019_/Q hold945/A _13827_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11120_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08303__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 hold870/A vssd1 vssd1 vccd1 vccd1 hold870/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 hold881/A vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11051_/X sky130_fd_sc_hd__or2_1
Xhold892 hold892/A vssd1 vssd1 vccd1 vccd1 hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ _09999_/Y _10000_/X _10002_/C _14961_/Q vssd1 vssd1 vccd1 vccd1 _10003_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__10271__C _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2260 _11664_/X vssd1 vssd1 vccd1 vccd1 _14467_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2271 _14016_/Q vssd1 vssd1 vccd1 vccd1 hold2271/X sky130_fd_sc_hd__dlygate4sd3_1
X_14810_ _15246_/CLK hold288/X vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2282 _07425_/X vssd1 vssd1 vccd1 vccd1 _14055_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07119__A0 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12338__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2293 _14144_/Q vssd1 vssd1 vccd1 vccd1 hold2293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1570 _07027_/X vssd1 vssd1 vccd1 vccd1 _13844_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1581 _14797_/Q vssd1 vssd1 vccd1 vccd1 hold1581/X sky130_fd_sc_hd__dlygate4sd3_1
X_14741_ _15382_/CLK _14741_/D vssd1 vssd1 vccd1 vccd1 _14741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _13708_/A1 hold2247/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11953_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12663__A1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1592 _07082_/X vssd1 vssd1 vccd1 vccd1 _13895_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _10717_/B _10719_/C _11091_/A _10903_/Y vssd1 vssd1 vccd1 vccd1 _11091_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _15377_/CLK hold722/X vssd1 vssd1 vccd1 vccd1 hold721/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ hold1243/X _13705_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13623_ input37/X _13636_/B vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__or2_1
Xclkbuf_2_3_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_10835_ _10835_/A _10835_/B vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13090__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15428_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13554_ _13554_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__or2_1
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10766_ hold735/A hold903/A hold309/A hold759/A _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _10767_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _12327_/A _12504_/X _12502_/X vssd1 vssd1 vccd1 vccd1 _13147_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_129_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__C _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ _11620_/A _11378_/C _10469_/X _10468_/X _11537_/B vssd1 vssd1 vccd1 vccd1
+ _10702_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13485_ _13492_/A hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__and2_1
XFILLER_0_125_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15224_ _15226_/CLK _15224_/D vssd1 vssd1 vccd1 vccd1 _15224_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_152_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12436_ _12642_/A1 _12435_/X _12700_/S0 vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15155_ _15316_/CLK _15155_/D vssd1 vssd1 vccd1 vccd1 _15155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12434__S _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ hold859/A _13800_/Q _12566_/S vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10743__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07528__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ _15390_/CLK hold986/X vssd1 vssd1 vccd1 vccd1 hold985/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _11499_/B1 _11311_/Y _11313_/Y _11315_/Y _11317_/Y vssd1 vssd1 vccd1 vccd1
+ _11318_/X sky130_fd_sc_hd__o32a_1
X_12298_ _15349_/Q _11729_/B _12296_/X _12297_/X _11997_/A vssd1 vssd1 vccd1 vccd1
+ _12301_/B sky130_fd_sc_hd__a2111o_1
X_15086_ _15375_/CLK hold348/X vssd1 vssd1 vccd1 vccd1 hold347/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14037_ _14083_/CLK _14037_/D vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
X_11249_ _11248_/B _11348_/B _11248_/A vssd1 vssd1 vccd1 vccd1 _11250_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11154__A1 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14939_ _15389_/CLK _14939_/D vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12654__A1 _13387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__B1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _14581_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08460_ _12247_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08460_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09979__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07411_ _13501_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _14041_/D sky130_fd_sc_hd__and2_1
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08391_ _08306_/A _08306_/B _08306_/C vssd1 vssd1 vccd1 vccd1 _08393_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09698__B _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__S _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15320_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11513__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07342_ _14057_/Q _07885_/A vssd1 vssd1 vccd1 vccd1 _07342_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09283__B1 _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10968__A1 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2752_A _10918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ _15222_/Q _14966_/Q vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09012_ _09253_/A _09712_/B _09011_/C _09011_/D vssd1 vssd1 vccd1 vccd1 _09012_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10356__C _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__A2_N _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12395__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__A0 _15058_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12344__S _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08123__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09914_ _09914_/A _09914_/B _09914_/C vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__nand3_1
Xfanout602 _09860_/B vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__clkbuf_4
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 _10022_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__buf_6
Xfanout624 _10033_/A vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout635 _15201_/Q vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout646 _08892_/A vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__buf_4
X_09845_ _09846_/B _14961_/Q _10108_/C _10000_/A vssd1 vssd1 vccd1 vccd1 _09847_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout657 _15067_/Q vssd1 vssd1 vccd1 vccd1 _13681_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 _13708_/A1 vssd1 vssd1 vccd1 vccd1 _13741_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout570_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__A1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 hold2735/X vssd1 vssd1 vccd1 vccd1 _13704_/A1 sky130_fd_sc_hd__buf_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout668_A _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09491_/A _09488_/Y _09628_/A _09775_/X _09626_/A vssd1 vssd1 vccd1 vccd1
+ _09776_/X sky130_fd_sc_hd__o311a_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ _13512_/A0 hold1207/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06988_/X sky130_fd_sc_hd__mux2_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07173__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08727_ _08593_/X _08596_/X _08725_/X _08726_/Y vssd1 vssd1 vccd1 vccd1 _08727_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13020__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout835_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08313__A2 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08869_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08658_/Y sky130_fd_sc_hd__nor2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08793__A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _13715_/A1 hold1465/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07609_/X sky130_fd_sc_hd__mux2_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08589_ _08589_/A _08589_/B _08589_/C vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__and3_1
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10620_ _10620_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__and2_1
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10551_ _10547_/Y _10549_/X _10337_/Y _10380_/X vssd1 vssd1 vccd1 vccd1 _10553_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07824__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13270_ input160/X fanout6/X fanout4/X input128/X vssd1 vssd1 vccd1 vccd1 _13270_/X
+ sky130_fd_sc_hd__a22o_1
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10482_/Y sky130_fd_sc_hd__xnor2_2
X_12221_ _12221_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12581__B1 _13150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _14887_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__or2_1
XANTENNA__11378__B _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11103_ _11288_/A1 _11102_/Y _10950_/X vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12083_ hold2435/X _12099_/A2 _12082_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12083_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11136__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11034_ _11033_/A _11033_/B _11033_/C _11033_/D vssd1 vssd1 vccd1 vccd1 _11035_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08001__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13085__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2090 _07137_/X vssd1 vssd1 vccd1 vccd1 _13947_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07083__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ hold1773/X hold2233/X _12991_/S vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__mux2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08304__A2 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _15365_/CLK _14724_/D vssd1 vssd1 vccd1 vccd1 _14724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _13691_/A1 hold1795/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__A2 _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _15435_/CLK hold454/X vssd1 vssd1 vccd1 vccd1 hold453/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ hold671/X _13655_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold672/A sky130_fd_sc_hd__mux2_1
XFILLER_0_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13606_ _07426_/A _13625_/C _13605_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15330_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13597__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08068__A1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ _10817_/B _10817_/C _10817_/A vssd1 vssd1 vccd1 vccd1 _10819_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13061__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14586_ _15458_/CLK hold266/X vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__dfxtp_1
X_11798_ hold1955/X _13652_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13537_ hold2354/X _13797_/A2 _13536_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15294_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10749_ _11108_/B _10749_/B vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13468_ _13468_/A _13468_/B vssd1 vssd1 vccd1 vccd1 _13468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11569__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15207_ _15226_/CLK _15207_/D vssd1 vssd1 vccd1 vccd1 _15207_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_211_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12419_ _12644_/A1 _12414_/X _12418_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12420_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10473__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput205 _14188_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[18] sky130_fd_sc_hd__buf_12
X_13399_ _13404_/A _13399_/B vssd1 vssd1 vccd1 vccd1 _15190_/D sky130_fd_sc_hd__and2_1
XFILLER_0_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput216 _14198_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[28] sky130_fd_sc_hd__buf_12
XFILLER_0_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput227 _14179_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[9] sky130_fd_sc_hd__buf_12
XFILLER_0_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15138_ _15299_/CLK _15138_/D vssd1 vssd1 vccd1 vccd1 _15138_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput238 _14443_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[19] sky130_fd_sc_hd__buf_12
Xoutput249 _14453_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[29] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09981__B _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _10873_/A _08012_/B vssd1 vssd1 vccd1 vccd1 _07961_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15069_ _15261_/CLK _15069_/D vssd1 vssd1 vccd1 vccd1 _15069_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_4_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15299_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_208_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06911_ _15342_/Q vssd1 vssd1 vccd1 vccd1 _07862_/B sky130_fd_sc_hd__inv_2
X_07891_ _10873_/A _08075_/B _07890_/C _07958_/A vssd1 vssd1 vccd1 vccd1 _07894_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10920__B _13460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09630_ _09918_/A _13444_/B _13361_/B _08256_/A _09629_/Y vssd1 vssd1 vccd1 vccd1
+ _09630_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09561_ _10002_/C _10010_/B vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13723__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ _08512_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _08514_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10638__B1 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12722__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _15151_/Q _09925_/A2 _07390_/A vssd1 vssd1 vccd1 vccd1 _09492_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07721__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08443_ _08542_/A _08544_/C vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__and2_1
XFILLER_0_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08374_ _12252_/B _08374_/B vssd1 vssd1 vccd1 vccd1 _08374_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ _11286_/A _09341_/A _08530_/B _09481_/A vssd1 vssd1 vccd1 vccd1 _07326_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_A _13716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _11168_/A _10304_/C vssd1 vssd1 vccd1 vccd1 _08846_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ hold1153/X _13655_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07187_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07168__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout785_A _14942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout410 _07115_/Y vssd1 vssd1 vccd1 vccd1 _07147_/S sky130_fd_sc_hd__clkbuf_16
Xfanout421 _13204_/Y vssd1 vssd1 vccd1 vccd1 _13220_/S sky130_fd_sc_hd__clkbuf_16
Xfanout432 _11763_/Y vssd1 vssd1 vccd1 vccd1 _11795_/S sky130_fd_sc_hd__clkbuf_16
Xfanout443 _13591_/A2 vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__buf_4
Xfanout454 _07981_/A vssd1 vssd1 vccd1 vccd1 _13636_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__10830__B _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _12129_/A2 vssd1 vssd1 vccd1 vccd1 _12099_/A2 sky130_fd_sc_hd__buf_4
Xfanout476 _07359_/X vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__buf_4
X_09828_ _10185_/A _10830_/B _09828_/C _09828_/D vssd1 vssd1 vccd1 vccd1 _09828_/X
+ sky130_fd_sc_hd__and4_1
Xfanout487 _12124_/D vssd1 vssd1 vccd1 vccd1 _12131_/B sky130_fd_sc_hd__clkbuf_4
Xfanout498 _06943_/Y vssd1 vssd1 vccd1 vccd1 _12844_/A1 sky130_fd_sc_hd__buf_8
XFILLER_0_198_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09759_ _09760_/A _09475_/B _09760_/B _09759_/D vssd1 vssd1 vccd1 vccd1 _09759_/X
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__12618__A1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A1 input136/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ _12770_/A _12770_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__or3b_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07631__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ hold1911/X _13741_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 _11721_/X sky130_fd_sc_hd__mux2_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _15313_/CLK _14440_/D vssd1 vssd1 vccd1 vccd1 _14440_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09247__B1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13043__A1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11652_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_182_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _10519_/A _10519_/B _10521_/X vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14371_ _15270_/CLK _14371_/D vssd1 vssd1 vccd1 vccd1 _14371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13322_ input83/X fanout2/X _13321_/X vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08470__A1 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ _10534_/A _10534_/B _10534_/C vssd1 vssd1 vccd1 vccd1 _10534_/X sky130_fd_sc_hd__and3_2
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13588__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08470__B2 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11389__A _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13253_ input90/X fanout1/X _13252_/X vssd1 vssd1 vccd1 vccd1 _13254_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ _10464_/B _10464_/C _10464_/A vssd1 vssd1 vccd1 vccd1 _10467_/C sky130_fd_sc_hd__o21ai_1
X_12204_ hold917/A _15261_/Q _12237_/S vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__mux2_1
X_10396_ _10395_/B _10736_/A vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_103_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13184_ _13393_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _15049_/D sky130_fd_sc_hd__and2_1
XANTENNA__10565__C1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output168_A _15180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08773__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12135_ _12068_/A _12195_/A2 _12134_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12135_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07806__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ _12066_/A _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12066_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09722__A1 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__B2 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _11570_/A _11409_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11201_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12013__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__B _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13282__A1 input133/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__B1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ _13068_/A1 _12965_/X _12967_/X vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06946__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07541__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _15449_/CLK hold492/X vssd1 vssd1 vccd1 vccd1 hold491/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ _13674_/A1 hold2129/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10468__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _13885_/Q hold839/A hold685/A hold867/A _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12899_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _15278_/CLK hold352/X vssd1 vssd1 vccd1 vccd1 hold351/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09789__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14569_ _14569_/CLK hold248/X vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07110_ _15066_/Q hold1807/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07110_/X sky130_fd_sc_hd__mux2_1
X_08090_ _08677_/A _11517_/A _08089_/C _08161_/B vssd1 vssd1 vccd1 vccd1 _08093_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07041_ hold1139/X _13679_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 _07041_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08213__A1 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold2715_A _11102_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13718__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _08992_/A1 _08985_/Y _08987_/Y _08989_/Y _08991_/Y vssd1 vssd1 vccd1 vccd1
+ _08992_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07716__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2804 _12339_/X vssd1 vssd1 vccd1 vccd1 hold2804/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2815 _14659_/Q vssd1 vssd1 vccd1 vccd1 hold2815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2826 _15334_/Q vssd1 vssd1 vccd1 vccd1 hold2826/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07943_ _15393_/Q _14528_/Q hold719/A _14752_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07943_/X sky130_fd_sc_hd__mux4_1
Xhold2837 _15338_/Q vssd1 vssd1 vccd1 vccd1 hold2837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2848 _15330_/Q vssd1 vssd1 vccd1 vccd1 hold2848/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09713__A1 _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2859 _15341_/Q vssd1 vssd1 vccd1 vccd1 hold2859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07874_ _15344_/Q _11729_/B _07872_/X _07873_/X _11997_/A vssd1 vssd1 vccd1 vccd1
+ _07878_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09613_ _09471_/B _09470_/Y _09610_/Y _09611_/X vssd1 vssd1 vccd1 vccd1 _09759_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09544_ _10700_/A _09676_/D _09543_/C _09673_/A vssd1 vssd1 vccd1 vccd1 _09545_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13273__A1 input130/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09232__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ _09760_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_A _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08426_ _08519_/B _08427_/B _08427_/C vssd1 vssd1 vccd1 vccd1 _08524_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08357_ _08877_/A _08356_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08357_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08790__B _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09378__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07308_ _08244_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07324_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08288_ _10873_/A _09437_/A _08234_/A _08232_/A vssd1 vssd1 vccd1 vccd1 _08329_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07239_ _15226_/Q _14970_/Q vssd1 vssd1 vccd1 vccd1 _07240_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13201__B _13201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12536__B1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ _10426_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10250_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08204__A1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _10020_/A _10020_/B _10028_/B _10026_/X vssd1 vssd1 vccd1 vccd1 _10191_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07626__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _15191_/CLK _13940_/D vssd1 vssd1 vccd1 vccd1 _13940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11511__A1 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _15270_/CLK _13871_/D vssd1 vssd1 vccd1 vccd1 _13871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12822_ _14801_/Q _14513_/Q hold615/A _14737_/Q _12915_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12822_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13264__A1 input158/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12698__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08366__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12753_ _13668_/A1 _13103_/A2 _13078_/B1 _13189_/B vssd1 vssd1 vccd1 vccd1 _12753_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11704_ hold2023/X _13724_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11704_/X sky130_fd_sc_hd__mux2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12684_ hold881/A _13909_/Q _12735_/S vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14909_/CLK hold490/X vssd1 vssd1 vccd1 vccd1 hold489/A sky130_fd_sc_hd__dfxtp_1
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11636_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14354_ _15093_/CLK _14354_/D vssd1 vssd1 vccd1 vccd1 _14354_/Q sky130_fd_sc_hd__dfxtp_1
X_11566_ _11566_/A _15226_/Q vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13305_ _13317_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _15121_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10517_ _10517_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14285_ _15446_/CLK _14285_/D vssd1 vssd1 vccd1 vccd1 _14285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ hold535/X _13748_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold536/A sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ _11596_/A _11597_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _10450_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12622__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13167_ _13168_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _15032_/D sky130_fd_sc_hd__nor2_1
X_10379_ _10380_/A _10380_/B _10439_/B _10380_/D vssd1 vssd1 vccd1 vccd1 _10379_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__09962__D _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _14999_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12118_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11566__B _15226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ hold227/A _14329_/Q hold557/A _13989_/Q _13091_/S _13098_/S1 vssd1 vssd1
+ vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09036__B _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12049_ _12063_/A _12049_/B vssd1 vssd1 vccd1 vccd1 _14837_/D sky130_fd_sc_hd__and2_1
XANTENNA__12925__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07590_ hold2822/X hold1933/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07590_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13255__A1 input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12689__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12463__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08131__B1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07336__A_N _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ _09260_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08211_ _08893_/A _08809_/B _08809_/D _08901_/A vssd1 vssd1 vccd1 vccd1 _08212_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09191_ _09190_/B _09190_/C _09190_/A vssd1 vssd1 vccd1 vccd1 _09191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13302__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08142_ _09008_/A _08776_/A _10507_/A _11550_/A vssd1 vssd1 vccd1 vccd1 _08144_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10645__B _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07300__A _15219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10241__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ _08312_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ hold687/X _13662_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 hold688/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2601 _15343_/Q vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_80_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11476__B _13466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2612 _14449_/Q vssd1 vssd1 vccd1 vccd1 _06914_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08975_ hold249/A _14313_/Q _14604_/Q _13973_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08975_/X sky130_fd_sc_hd__mux4_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _07862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2623 _15296_/Q vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__buf_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2634 _14980_/Q vssd1 vssd1 vccd1 vccd1 hold2634/X sky130_fd_sc_hd__buf_2
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1900 _07161_/X vssd1 vssd1 vccd1 vccd1 _13969_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2645 _08861_/X vssd1 vssd1 vccd1 vccd1 _14437_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2656 _14824_/Q vssd1 vssd1 vccd1 vccd1 hold2656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1911 _14517_/Q vssd1 vssd1 vccd1 vccd1 hold1911/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _07926_/A _07926_/B vssd1 vssd1 vccd1 vccd1 _07926_/Y sky130_fd_sc_hd__nand2_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2667 _14819_/Q vssd1 vssd1 vccd1 vccd1 hold2667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1922 _07509_/X vssd1 vssd1 vccd1 vccd1 _14137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1933 _14214_/Q vssd1 vssd1 vccd1 vccd1 hold1933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2678 _14830_/Q vssd1 vssd1 vccd1 vccd1 hold2678/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2689 _08186_/X vssd1 vssd1 vccd1 vccd1 _14430_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07970__A _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1944 _07151_/X vssd1 vssd1 vccd1 vccd1 _13959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1955 _14622_/Q vssd1 vssd1 vccd1 vccd1 hold1955/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ hold195/A hold95/A _07857_/C _07857_/D vssd1 vssd1 vccd1 vccd1 _07857_/X
+ sky130_fd_sc_hd__or4_1
Xhold1966 _07139_/X vssd1 vssd1 vccd1 vccd1 _13949_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1977 _14387_/Q vssd1 vssd1 vccd1 vccd1 hold1977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1988 _07769_/X vssd1 vssd1 vccd1 vccd1 _14385_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1999 _13847_/Q vssd1 vssd1 vccd1 vccd1 hold1999/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13246__A1 input140/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07788_ hold925/X _13693_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold926/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07181__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09527_ _09527_/A _09527_/B _09527_/C vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09457_/A _09587_/A _09557_/A _09457_/D vssd1 vssd1 vccd1 vccd1 _09459_/C
+ sky130_fd_sc_hd__o22ai_4
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _08473_/A _08300_/B _08503_/A vssd1 vssd1 vccd1 vccd1 _08410_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__13549__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _09285_/A _09285_/B _09285_/C vssd1 vssd1 vccd1 vccd1 _09390_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _11420_/A _11551_/B _11420_/C vssd1 vssd1 vccd1 vccd1 _11420_/X sky130_fd_sc_hd__and3_1
XFILLER_0_163_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _11541_/A _11351_/B _11620_/B _15221_/Q vssd1 vssd1 vccd1 vccd1 _11352_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08025__B _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _11168_/A _10304_/C _10304_/D _11605_/A vssd1 vssd1 vccd1 vccd1 _10306_/C
+ sky130_fd_sc_hd__a22o_1
X_14070_ _15225_/CLK _14070_/D vssd1 vssd1 vccd1 vccd1 _14070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _11282_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08189__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ hold1601/X hold963/X hold411/X hold1535/X _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13021_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10233_ _10233_/A _10409_/B _10233_/C vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__or3_1
XANTENNA__09137__A _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _10164_/A _10336_/A _10164_/C vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__or3_2
XANTENNA__10091__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__A _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ _14353_/Q _14257_/Q hold841/A _14129_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10096_/B sky130_fd_sc_hd__mux4_1
X_14972_ _14972_/CLK _14972_/D vssd1 vssd1 vccd1 vccd1 _14972_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10299__A1 _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13923_ _15456_/CLK _13923_/D vssd1 vssd1 vccd1 vccd1 _13923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08695__B _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13854_ _15093_/CLK _13854_/D vssd1 vssd1 vccd1 vccd1 _13854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07091__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _13080_/A1 _12804_/X _12802_/X vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13788__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13785_ hold265/X vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10997_ _10996_/A _10996_/B _10996_/C _10996_/D vssd1 vssd1 vccd1 vccd1 _10997_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12917_/A1 _12735_/X _12844_/A1 vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__a21o_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08664__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10168__D _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15455_ _15455_/CLK hold576/X vssd1 vssd1 vccd1 vccd1 hold575/A sky130_fd_sc_hd__dfxtp_1
X_12667_ _12692_/A1 _12666_/X _12366_/A vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13096__S0 _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ _15372_/CLK _14406_/D vssd1 vssd1 vccd1 vccd1 _14406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _11618_/A _11618_/B vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15386_ _15421_/CLK _15386_/D vssd1 vssd1 vccd1 vccd1 _15386_/Q sky130_fd_sc_hd__dfxtp_1
X_12598_ hold253/A hold817/A _14600_/Q _13969_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12598_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ _15080_/CLK hold852/X vssd1 vssd1 vccd1 vccd1 hold851/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11549_ _11402_/A _11401_/A _11401_/B _11403_/Y vssd1 vssd1 vccd1 vccd1 _11553_/A
+ sky130_fd_sc_hd__o31ai_1
Xhold507 hold507/A vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 hold518/A vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold529 hold529/A vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ _15222_/CLK _14268_/D vssd1 vssd1 vccd1 vccd1 _14268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09916__A1 _11287_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__A _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13219_ hold1541/X _13665_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08275__S0 _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _15087_/CLK _14199_/D vssd1 vssd1 vccd1 vccd1 _14199_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07927__B1 _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2413_A _15036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1207 _13807_/Q vssd1 vssd1 vccd1 vccd1 hold1207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _08760_/A _08760_/B vssd1 vssd1 vccd1 vccd1 _08760_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_139_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1218 _11958_/X vssd1 vssd1 vccd1 vccd1 _14778_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1229 _14328_/Q vssd1 vssd1 vccd1 vccd1 hold1229/X sky130_fd_sc_hd__dlygate4sd3_1
X_07711_ hold1263/X _12329_/A _07726_/S vssd1 vssd1 vccd1 vccd1 _07711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08691_ _08691_/A _08691_/B vssd1 vssd1 vccd1 vccd1 _08692_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07642_ hold1791/X _13748_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07642_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2782_A _14492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ _13404_/A _07573_/B vssd1 vssd1 vccd1 vccd1 _14198_/D sky130_fd_sc_hd__and2_1
XFILLER_0_177_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13731__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ _09309_/Y _09310_/X _09178_/Y _09180_/X vssd1 vssd1 vccd1 vccd1 _09314_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09510__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ _11320_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09243_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12347__S _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__A _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _09297_/B _09173_/C _09173_/A vssd1 vssd1 vccd1 vccd1 _09175_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11411__B1 _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _08869_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _08125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09080__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08056_ _14786_/Q hold789/A _14626_/Q _14722_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08057_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07007_ _13679_/A1 hold1953/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07007_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08266__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10822__C _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12911__B1 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput105 in1[17] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__clkbuf_1
Xinput116 in1[27] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_1
Xhold2420 _14858_/Q vssd1 vssd1 vccd1 vccd1 hold2420/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout865_A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput127 in1[8] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2431 _13573_/X vssd1 vssd1 vccd1 vccd1 _15312_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 in2[18] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__clkbuf_2
X_08958_ _09119_/A _08957_/B _08957_/Y _11473_/A vssd1 vssd1 vccd1 vccd1 _08958_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2442 _11474_/X vssd1 vssd1 vccd1 vccd1 _13404_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12810__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput149 in2[28] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_192_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2453 _12075_/X vssd1 vssd1 vccd1 vccd1 _14849_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2464 _13429_/X vssd1 vssd1 vccd1 vccd1 _15208_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2475 _14865_/Q vssd1 vssd1 vccd1 vccd1 hold2475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 _07091_/X vssd1 vssd1 vccd1 vccd1 _13904_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ _09344_/B _07910_/B vssd1 vssd1 vccd1 vccd1 _08637_/B sky130_fd_sc_hd__nor2_2
Xhold2486 _12187_/X vssd1 vssd1 vccd1 vccd1 _14904_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1741 _13955_/Q vssd1 vssd1 vccd1 vccd1 hold1741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1752 _07050_/X vssd1 vssd1 vccd1 vccd1 _13866_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08889_ _09858_/A _08888_/X _08887_/X vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__a21bo_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2497 _15351_/Q vssd1 vssd1 vccd1 vccd1 _08107_/A sky130_fd_sc_hd__clkbuf_4
Xhold1763 _14476_/Q vssd1 vssd1 vccd1 vccd1 hold1763/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1774 _11857_/X vssd1 vssd1 vccd1 vccd1 _14680_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1785 _14533_/Q vssd1 vssd1 vccd1 vccd1 hold1785/X sky130_fd_sc_hd__dlygate4sd3_1
X_10920_ _13749_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _10920_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09404__B _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1796 _11936_/X vssd1 vssd1 vccd1 vccd1 _14756_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10851_ _10850_/B _10850_/C _10850_/A vssd1 vssd1 vccd1 vccd1 _10851_/Y sky130_fd_sc_hd__a21oi_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12978__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_160_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _14441_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13570_/X sky130_fd_sc_hd__or2_1
X_10782_ _10782_/A _10970_/A vssd1 vssd1 vccd1 vccd1 _10792_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10453__A1 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _15366_/Q _15269_/Q hold527/A hold457/A _12560_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12521_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clk_A clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15243_/CLK _15240_/D vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12452_ _13027_/A _12452_/B _12452_/C vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__and3_1
XFILLER_0_136_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12825__S0 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11403_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11403_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_leaf_175_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15171_ _15365_/CLK _15171_/D vssd1 vssd1 vccd1 vccd1 _15171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12383_ _15393_/Q _14528_/Q hold719/A _14752_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12383_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10756__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ _14472_/CLK _14122_/D vssd1 vssd1 vccd1 vccd1 _14122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11334_ _11334_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11336_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13596__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ _15422_/CLK _14053_/D vssd1 vssd1 vccd1 vccd1 hold313/A sky130_fd_sc_hd__dfxtp_1
X_11265_ _11460_/A _11264_/B _11328_/B _11264_/D vssd1 vssd1 vccd1 vccd1 _11265_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10508__A2 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07086__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _10918_/X _13104_/A2 _13003_/X vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__a21o_1
X_10216_ _10392_/B _10215_/X _10065_/B _10065_/Y vssd1 vssd1 vccd1 vccd1 _10263_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11196_ _11564_/A _11378_/D _11196_/C _11382_/A vssd1 vssd1 vccd1 vccd1 _11382_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10147_ _10312_/B _10145_/X _10007_/X _10011_/B vssd1 vssd1 vccd1 vccd1 _10148_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13458__A1 _12286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07814__S _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14955_ _14955_/CLK _14955_/D vssd1 vssd1 vccd1 vccd1 _14955_/Q sky130_fd_sc_hd__dfxtp_1
X_10078_ _07261_/A _07319_/D _09915_/X _10077_/Y vssd1 vssd1 vccd1 vccd1 _10078_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13906_ _15439_/CLK _13906_/D vssd1 vssd1 vccd1 vccd1 _13906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08885__A1 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14886_ _14989_/CLK _14886_/D vssd1 vssd1 vccd1 vccd1 _14886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12681__A2 _13154_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09509__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13837_ _15264_/CLK _13837_/D vssd1 vssd1 vccd1 vccd1 _13837_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08980__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11316__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_128_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13768_ hold247/X vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12719_ _12844_/A1 _12714_/X _12718_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12720_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__10476__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ hold609/X _13732_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold610/A sky130_fd_sc_hd__mux2_1
XFILLER_0_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15438_ _15438_/CLK _15438_/D vssd1 vssd1 vccd1 vccd1 _15438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15369_ _15369_/CLK hold472/X vssd1 vssd1 vccd1 vccd1 hold471/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10747__A2 _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold315 hold315/A vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold337 hold337/A vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold348 hold348/A vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ _09930_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _09932_/C sky130_fd_sc_hd__or2_1
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold359 hold359/A vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold2628_A _14977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10642__C _14954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout806 _12365_/S1 vssd1 vssd1 vccd1 vccd1 _12668_/A1 sky130_fd_sc_hd__clkbuf_8
X_09861_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout817 _13098_/S1 vssd1 vssd1 vccd1 vccd1 _13099_/S1 sky130_fd_sc_hd__clkbuf_8
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout828 _12365_/S0 vssd1 vssd1 vccd1 vccd1 _12560_/S sky130_fd_sc_hd__buf_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08573__B1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__B2 _15345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _12991_/S sky130_fd_sc_hd__clkbuf_4
X_08812_ _08812_/A _08922_/B _08812_/C vssd1 vssd1 vccd1 vccd1 _08814_/B sky130_fd_sc_hd__nand3_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13726__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _10244_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__or2_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _07514_/X vssd1 vssd1 vccd1 vccd1 _14139_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 _14699_/Q vssd1 vssd1 vccd1 vccd1 hold1015/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _07018_/X vssd1 vssd1 vccd1 vccd1 _13835_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07724__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08743_ _08743_/A _09346_/B _08743_/C vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__or3_1
Xhold1037 _14712_/Q vssd1 vssd1 vccd1 vccd1 hold1037/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 _13723_/X vssd1 vssd1 vccd1 vccd1 _15433_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1059 _14670_/Q vssd1 vssd1 vccd1 vccd1 hold1059/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13027__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _08674_/A _08674_/B vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ hold1925/X _13698_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07556_ _13393_/A hold135/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__and2_1
XANTENNA__09825__B1 _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__B2 _13197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout613_A _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ hold1453/X _13693_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07487_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10986__A2 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09226_ _09514_/A _09225_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_9_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ _09157_/A _09157_/B _09157_/C vssd1 vssd1 vccd1 vccd1 _09159_/A sky130_fd_sc_hd__and3_1
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ _08106_/Y _08108_/B vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_142_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _14438_/Q _09087_/C _09087_/A vssd1 vssd1 vccd1 vccd1 _09089_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__and2_1
XFILLER_0_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12106__A _14993_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 hold860/A vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08303__B _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 hold871/A vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 hold882/A vssd1 vssd1 vccd1 vccd1 hold882/X sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _10868_/B _10870_/B _10868_/A vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__o21ba_1
Xhold893 hold893/A vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10001_ _10002_/C _14961_/Q _09999_/Y _10000_/X vssd1 vssd1 vccd1 vccd1 _10003_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12540__S _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2250 _07108_/X vssd1 vssd1 vccd1 vccd1 _13921_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2261 _15264_/Q vssd1 vssd1 vccd1 vccd1 hold2261/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07634__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2272 _07209_/X vssd1 vssd1 vccd1 vccd1 _14016_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2283 _14916_/Q vssd1 vssd1 vccd1 vccd1 _13477_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2294 _07519_/X vssd1 vssd1 vccd1 vccd1 _14144_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1560 _07651_/X vssd1 vssd1 vccd1 vccd1 _14272_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _15408_/CLK _14740_/D vssd1 vssd1 vccd1 vccd1 _14740_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1571 _13952_/Q vssd1 vssd1 vccd1 vccd1 hold1571/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ _15060_/Q hold1715/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__mux2_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1582 _11978_/X vssd1 vssd1 vccd1 vccd1 _14797_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1593 _14375_/Q vssd1 vssd1 vccd1 vccd1 hold1593/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _11085_/B _10901_/Y _10675_/Y _10719_/X vssd1 vssd1 vccd1 vccd1 _10903_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _15408_/CLK _14671_/D vssd1 vssd1 vccd1 vccd1 _14671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ hold933/X _13704_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold934/A sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12776__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ _08741_/A _13625_/C _13621_/X _13622_/C1 vssd1 vssd1 vccd1 vccd1 _15338_/D
+ sky130_fd_sc_hd__o211a_1
X_10834_ _10832_/X _10834_/B vssd1 vssd1 vccd1 vccd1 _10835_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_211_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ _08345_/B _13591_/A2 _13552_/X _13541_/A vssd1 vssd1 vccd1 vccd1 _13553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10765_ _11509_/A _10765_/B vssd1 vssd1 vccd1 vccd1 _10765_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _08248_/Y _12325_/B _12503_/X vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13484_ _13490_/A hold97/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__and2_1
XANTENNA__09300__D _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10696_ _10696_/A _10696_/B vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12179__A1 _12112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15223_ _15226_/CLK _15223_/D vssd1 vssd1 vccd1 vccd1 _15223_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12435_ hold435/A _13931_/Q _12441_/S vssd1 vssd1 vccd1 vccd1 _12435_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09044__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12715__S _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13400__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15154_ _15316_/CLK _15154_/D vssd1 vssd1 vccd1 vccd1 _15154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12366_ _12366_/A _12366_/B vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__or2_1
XFILLER_0_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14105_ _14105_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _14105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _11507_/A _11316_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _11317_/Y sky130_fd_sc_hd__o21ai_1
X_15085_ _15374_/CLK hold944/X vssd1 vssd1 vccd1 vccd1 hold943/A sky130_fd_sc_hd__dfxtp_1
X_12297_ _15348_/Q _07744_/A _14089_/Q _13240_/A vssd1 vssd1 vccd1 vccd1 _12297_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ _14083_/CLK _14036_/D vssd1 vssd1 vccd1 vccd1 _14036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11248_ _11248_/A _11248_/B _11348_/B vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__nand3_2
XANTENNA__11154__A2 _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__A1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11179_ _11179_/A _11179_/B _11179_/C vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__and3_1
XFILLER_0_59_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07544__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14938_ _14972_/CLK _14938_/D vssd1 vssd1 vccd1 vccd1 _14938_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12654__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09979__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ _14876_/CLK _14869_/D vssd1 vssd1 vccd1 vccd1 _14869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07410_ _13501_/A _07410_/B vssd1 vssd1 vccd1 vccd1 _14040_/D sky130_fd_sc_hd__and2_1
XANTENNA__11590__A _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ _08389_/B _08389_/C _08389_/A vssd1 vssd1 vccd1 vccd1 _08393_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08375__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09807__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__A1 _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07341_ _07852_/A _07341_/B _07408_/A _07407_/A vssd1 vssd1 vccd1 vccd1 _07885_/A
+ sky130_fd_sc_hd__or4b_4
XANTENNA__09283__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2578_A _14432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09283__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10637__C _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__A2 _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07272_ _15222_/Q _14966_/Q vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__or2_1
X_09011_ _09253_/A _09712_/B _09011_/C _09011_/D vssd1 vssd1 vccd1 vccd1 _09011_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10356__D _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2745_A _15174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07719__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _11474_/A2 _09911_/Y _09912_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__o211a_1
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _15210_/Q vssd1 vssd1 vccd1 vccd1 _09860_/B sky130_fd_sc_hd__buf_8
XFILLER_0_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout614 _10022_/A vssd1 vssd1 vccd1 vccd1 _11563_/A sky130_fd_sc_hd__clkbuf_8
Xfanout625 _10033_/A vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__buf_4
XANTENNA__08546__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_A _07677_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout636 _08012_/B vssd1 vssd1 vccd1 vccd1 _08776_/A sky130_fd_sc_hd__buf_4
X_09844_ _09841_/X _09842_/Y _09690_/B _09692_/B vssd1 vssd1 vccd1 vccd1 _09896_/B
+ sky130_fd_sc_hd__o211a_1
Xfanout647 _15198_/Q vssd1 vssd1 vccd1 vccd1 _08892_/A sky130_fd_sc_hd__clkbuf_8
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout658 _13746_/A1 vssd1 vssd1 vccd1 vccd1 _13680_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 _13708_/A1 vssd1 vssd1 vccd1 vccd1 _13675_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09775_/A _09775_/B _09626_/B vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__or3b_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ _13659_/A1 hold1935/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06987_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout563_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08726_ _08725_/A _08725_/B _08621_/B vssd1 vssd1 vccd1 vccd1 _08726_/Y sky130_fd_sc_hd__o21bai_2
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08657_ _14342_/Q _14246_/Q _14406_/Q _14118_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08658_/B sky130_fd_sc_hd__mux4_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout730_A _14958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08793__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11704__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _13714_/A1 hold823/X _07609_/S vssd1 vssd1 vccd1 vccd1 hold824/A sky130_fd_sc_hd__mux2_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _08480_/A _08480_/B _08480_/C vssd1 vssd1 vccd1 vccd1 _08589_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07539_ hold1599/X _13743_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 _07539_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ _10337_/Y _10380_/X _10547_/Y _10549_/X vssd1 vssd1 vccd1 vccd1 _10553_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _13390_/B vssd1 vssd1 vccd1 vccd1 _09209_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _10479_/X _10481_/B vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__S _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ hold2757/X _12254_/A _12256_/A vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12030__A0 hold2509/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12581__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ hold2607/X _12173_/A2 _12150_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11378__C _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _06941_/Y _12256_/A _10956_/Y _10957_/X _11101_/X vssd1 vssd1 vccd1 vccd1
+ _11102_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_0_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12082_ _14981_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12082_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_124_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold690 hold690/A vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12869__C1 _06944_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13530__A0 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12333__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11033_ _11033_/A _11033_/B _11033_/C _11033_/D vssd1 vssd1 vccd1 vccd1 _11035_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2080 _07166_/X vssd1 vssd1 vccd1 vccd1 _13974_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2091 _13880_/Q vssd1 vssd1 vccd1 vccd1 hold2091/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ hold715/X hold2249/X _12991_/S vssd1 vssd1 vccd1 vccd1 _12984_/X sky130_fd_sc_hd__mux2_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1390 _11960_/X vssd1 vssd1 vccd1 vccd1 _14780_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10647__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ _13657_/A1 hold1445/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__mux2_1
X_14723_ _15305_/CLK _14723_/D vssd1 vssd1 vccd1 vccd1 _14723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _15360_/CLK hold854/X vssd1 vssd1 vccd1 vccd1 hold853/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ hold719/X _13654_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold720/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ input59/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__or2_1
X_10817_ _10817_/A _10817_/B _10817_/C vssd1 vssd1 vccd1 vccd1 _10819_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_185_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09265__A1 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14585_ _15421_/CLK hold260/X vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ hold855/X _13651_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold856/A sky130_fd_sc_hd__mux2_1
XFILLER_0_184_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13536_ _13536_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__or2_1
XFILLER_0_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10748_ _11108_/A _11108_/C _11110_/A vssd1 vssd1 vccd1 vccd1 _10749_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_165_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ _11478_/B _13466_/A _13466_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 _13467_/X
+ sky130_fd_sc_hd__o211a_1
X_10679_ _11550_/A _15219_/Q _11620_/B _11526_/A vssd1 vssd1 vccd1 vccd1 _10681_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07539__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15206_ _15226_/CLK _15206_/D vssd1 vssd1 vccd1 vccd1 _15206_/Q sky130_fd_sc_hd__dfxtp_1
X_12418_ _12474_/S1 _12415_/X _12417_/X vssd1 vssd1 vccd1 vccd1 _12418_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11569__B _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ _13479_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _15189_/D sky130_fd_sc_hd__and2_2
XANTENNA__10473__B _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput206 _14189_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[19] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput217 _14199_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[29] sky130_fd_sc_hd__buf_12
XFILLER_0_65_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _15301_/CLK _15137_/D vssd1 vssd1 vccd1 vccd1 _15137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput228 _15459_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[0] sky130_fd_sc_hd__buf_12
XFILLER_0_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12349_ _12343_/A _12348_/X _12366_/A vssd1 vssd1 vccd1 vccd1 _12349_/X sky130_fd_sc_hd__a21o_1
Xoutput239 _15460_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[1] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _15068_/CLK _15068_/D vssd1 vssd1 vccd1 vccd1 _15068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06910_ _15343_/Q vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__inv_2
X_14019_ _15387_/CLK _14019_/D vssd1 vssd1 vccd1 vccd1 _14019_/Q sky130_fd_sc_hd__dfxtp_1
X_07890_ _10873_/A _08075_/B _07890_/C _07958_/A vssd1 vssd1 vccd1 vccd1 _07963_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_65_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15207__D _15207_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09560_ _09557_/X _09558_/Y _09417_/B _09418_/Y vssd1 vssd1 vccd1 vccd1 _09602_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08511_ _08511_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10638__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10638__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2695_A _15190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09491_ _09491_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _13360_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13305__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ _13554_/B _08440_/Y _08441_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _14433_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07303__A _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08373_ _08358_/Y _08363_/Y _08372_/X _12241_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08374_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07324_ _07324_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _07326_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_46_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08464__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07255_ _07253_/Y _07255_/B vssd1 vssd1 vccd1 vccd1 _10951_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout409_A _07115_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12012__A0 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10249__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ hold681/X _13654_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold682/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08134__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__A1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
Xfanout400 _07577_/Y vssd1 vssd1 vccd1 vccd1 _07609_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__11118__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 _07080_/Y vssd1 vssd1 vccd1 vccd1 _07096_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout778_A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _13204_/Y vssd1 vssd1 vccd1 vccd1 _13236_/S sky130_fd_sc_hd__buf_12
XFILLER_0_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout433 _07778_/Y vssd1 vssd1 vccd1 vccd1 _07794_/S sky130_fd_sc_hd__clkbuf_16
Xfanout444 _07389_/Y vssd1 vssd1 vccd1 vccd1 _13591_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07184__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 _07012_/Y vssd1 vssd1 vccd1 vccd1 _07028_/S sky130_fd_sc_hd__clkbuf_16
Xfanout466 _12065_/Y vssd1 vssd1 vccd1 vccd1 _12129_/A2 sky130_fd_sc_hd__buf_4
X_09827_ _10185_/A _10830_/B _09828_/C _09828_/D vssd1 vssd1 vccd1 vccd1 _09827_/Y
+ sky130_fd_sc_hd__a22oi_2
Xfanout477 _13081_/A1 vssd1 vssd1 vccd1 vccd1 _13106_/A1 sky130_fd_sc_hd__buf_4
Xfanout488 _12124_/D vssd1 vssd1 vccd1 vccd1 _12128_/D sky130_fd_sc_hd__clkbuf_4
Xfanout499 _06943_/Y vssd1 vssd1 vccd1 vccd1 _12950_/S0 sky130_fd_sc_hd__buf_4
XFILLER_0_198_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ _09910_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__nor2_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08709_ _08709_/A _08805_/B _08709_/C vssd1 vssd1 vccd1 vccd1 _08712_/B sky130_fd_sc_hd__nand3_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09689_ _09686_/X _09687_/Y _09549_/X _09551_/Y vssd1 vssd1 vccd1 vccd1 _09690_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ hold649/X _13674_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 hold650/A sky130_fd_sc_hd__mux2_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ _11650_/B hold2528/X _11650_/Y _13369_/A vssd1 vssd1 vccd1 vccd1 _14455_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09247__A1 _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__C _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09247__B2 _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ _10599_/X _10601_/X _10951_/B vssd1 vssd1 vccd1 vccd1 _10602_/X sky130_fd_sc_hd__a21o_1
X_14370_ _15077_/CLK hold458/X vssd1 vssd1 vccd1 vccd1 hold457/A sky130_fd_sc_hd__dfxtp_1
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ input147/X fanout5/X fanout3/X input115/X vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ _10532_/B _10532_/C _10532_/A vssd1 vssd1 vccd1 vccd1 _10534_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ input154/X fanout6/X fanout4/X input122/X vssd1 vssd1 vccd1 vccd1 _13252_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10464_ _10464_/A _10464_/B _10464_/C vssd1 vssd1 vccd1 vccd1 _10635_/A sky130_fd_sc_hd__or3_2
XANTENNA__11389__B _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12554__A1 _13383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12203_ _15069_/Q _14362_/Q _12237_/S vssd1 vssd1 vccd1 vccd1 _12203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13183_ _13386_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _15048_/D sky130_fd_sc_hd__and2_1
X_10395_ _10736_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10395_/Y sky130_fd_sc_hd__nand2b_1
X_12134_ _14878_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12065_ _12096_/B _12096_/C _12124_/D vssd1 vssd1 vccd1 vccd1 _12065_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07094__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ _11409_/A _11537_/A _11623_/B _11570_/A vssd1 vssd1 vccd1 vccd1 _11018_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09722__A2 _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08210__C _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07822__S _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _13092_/A1 _12966_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__a21o_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14706_ _15411_/CLK _14706_/D vssd1 vssd1 vccd1 vccd1 _14706_/Q sky130_fd_sc_hd__dfxtp_1
X_11918_ _13673_/A1 hold2061/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11918_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13019__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08219__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ hold269/A hold335/A _14612_/Q _13981_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12898_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10468__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14637_ _15190_/CLK _14637_/D vssd1 vssd1 vccd1 vccd1 _14637_/Q sky130_fd_sc_hd__dfxtp_1
X_11849_ hold721/X _13736_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold722/A sky130_fd_sc_hd__mux2_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14568_ _15268_/CLK hold254/X vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12793__A1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13519_ _13519_/A0 hold1313/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13519_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2276_A _13472_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14499_ _15364_/CLK _14499_/D vssd1 vssd1 vccd1 vccd1 _14499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07040_ hold1687/X _13744_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08213__A2 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _08981_/A _08990_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08991_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_hold2610_A _15003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2805 _14155_/Q vssd1 vssd1 vccd1 vccd1 hold2805/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07942_ _08201_/A _07942_/B vssd1 vssd1 vccd1 vccd1 _07942_/Y sky130_fd_sc_hd__nor2_1
Xhold2816 _15038_/Q vssd1 vssd1 vccd1 vccd1 hold2816/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2827 _15337_/Q vssd1 vssd1 vccd1 vccd1 hold2827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2838 _15294_/Q vssd1 vssd1 vccd1 vccd1 hold2838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07955__A2_N _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2849 _15304_/Q vssd1 vssd1 vccd1 vccd1 hold2849/X sky130_fd_sc_hd__dlygate4sd3_1
X_07873_ _15342_/Q _07875_/B _14089_/Q _06909_/Y vssd1 vssd1 vccd1 vccd1 _07873_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09612_ _09610_/Y _09611_/X _09471_/B _09470_/Y vssd1 vssd1 vccd1 vccd1 _09760_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13734__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07732__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _10700_/A _09676_/D _09543_/C _09673_/A vssd1 vssd1 vccd1 vccd1 _09673_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_211_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09477__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout359_A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _09471_/X _09472_/Y _09328_/Y _09330_/Y vssd1 vssd1 vccd1 vccd1 _09475_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12481__B1 _13146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08425_ _08519_/B _08427_/B _08427_/C vssd1 vssd1 vccd1 vccd1 _08428_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_149_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout526_A _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08356_ _13871_/Q _13999_/Q _13839_/Q _13807_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08356_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07307_ _08702_/B _11541_/A vssd1 vssd1 vccd1 vccd1 _07308_/B sky130_fd_sc_hd__or2_1
XFILLER_0_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08287_ _13659_/A1 _12260_/A2 _12259_/A1 _13180_/B _08285_/Y vssd1 vssd1 vccd1 vccd1
+ _08287_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07179__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ _15226_/Q _14970_/Q vssd1 vssd1 vccd1 vccd1 _07240_/A sky130_fd_sc_hd__or2_1
XFILLER_0_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12536__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09401__A1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07169_ _13703_/A1 hold2001/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07169_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09401__B2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _10180_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12114__A _12114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13870_ _15077_/CLK _13870_/D vssd1 vssd1 vccd1 vccd1 _13870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07642__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ hold377/A _15281_/Q hold307/A _14382_/Q _12915_/S _12939_/S1 vssd1 vssd1
+ vccd1 vccd1 _12821_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12698__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10078__A2 _07319_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _13102_/A _12752_/B _12752_/C vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__and3_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ hold1841/X _13657_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__mux2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12683_ hold609/A _14540_/Q hold737/A _14764_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12683_/X sky130_fd_sc_hd__mux4_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14422_ _14485_/CLK _14422_/D vssd1 vssd1 vccd1 vccd1 _14422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13421__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _15196_/CLK _14353_/D vssd1 vssd1 vccd1 vccd1 _14353_/Q sky130_fd_sc_hd__dfxtp_1
X_11565_ _11565_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09640__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ input77/X fanout2/X _13303_/X vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07089__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10516_ _11340_/A _15221_/Q vssd1 vssd1 vccd1 vccd1 _10517_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14284_ _15411_/CLK hold674/X vssd1 vssd1 vccd1 vccd1 hold673/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output180_A _15191_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ hold469/A _13957_/Q hold361/A _13925_/Q _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _11497_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ hold451/X _13681_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold452/A sky130_fd_sc_hd__mux2_1
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10447_ _11596_/A _11597_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _10447_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_62_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12622__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ _13168_/A _13166_/B vssd1 vssd1 vccd1 vccd1 _15031_/D sky130_fd_sc_hd__nor2_1
X_10378_ _10439_/A _10376_/X _10196_/Y _10199_/Y vssd1 vssd1 vccd1 vccd1 _10380_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12117_ hold2461/X _12129_/A2 _12116_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12117_/X
+ sky130_fd_sc_hd__o211a_1
X_13097_ hold369/A hold385/A hold787/A hold991/A _13091_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13097_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_100_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12048_ _12114_/A hold2704/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12049_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12689__S1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ _15270_/CLK _13999_/D vssd1 vssd1 vccd1 vccd1 _13999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08131__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_190 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _08901_/A _08893_/A _08809_/B _08809_/D vssd1 vssd1 vccd1 vccd1 _08297_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_146_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11802__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09190_ _09190_/A _09190_/B _09190_/C vssd1 vssd1 vccd1 vccd1 _09324_/A sky130_fd_sc_hd__or3_2
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08141_ _11566_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__and2_1
XFILLER_0_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15220__D _15220_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07300__B _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ _13656_/A1 _12260_/A2 _12259_/A1 _13177_/B _08070_/Y vssd1 vssd1 vccd1 vccd1
+ _08072_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_109_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12518__A1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13729__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07023_ hold1089/X _13661_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07023_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07727__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07954__C _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__A1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08974_ _13570_/B _08972_/Y _08973_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _08974_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2602 _14981_/Q vssd1 vssd1 vccd1 vccd1 hold2602/X sky130_fd_sc_hd__buf_2
Xhold2613 _10576_/X vssd1 vssd1 vccd1 vccd1 _14449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2624 _13540_/X vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2635 _12147_/X vssd1 vssd1 vccd1 vccd1 _14884_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1901 _13967_/Q vssd1 vssd1 vccd1 vccd1 hold1901/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ hold2580/X _07812_/A _11104_/A _12262_/B _07922_/Y vssd1 vssd1 vccd1 vccd1
+ _07925_/X sky130_fd_sc_hd__a221o_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2646 _15166_/Q vssd1 vssd1 vccd1 vccd1 hold2646/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2657 _12022_/X vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1912 _11721_/X vssd1 vssd1 vccd1 vccd1 _14517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2668 _14816_/Q vssd1 vssd1 vccd1 vccd1 hold2668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1923 _14541_/Q vssd1 vssd1 vccd1 vccd1 hold1923/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2679 _12034_/X vssd1 vssd1 vccd1 vccd1 _12035_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1934 _07590_/X vssd1 vssd1 vccd1 vccd1 _14214_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07970__B _13412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1945 _14783_/Q vssd1 vssd1 vccd1 vccd1 hold1945/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ hold197/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07857_/D sky130_fd_sc_hd__nand2_1
Xhold1956 _11798_/X vssd1 vssd1 vccd1 vccd1 _14622_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10167__A2_N _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1967 _14389_/Q vssd1 vssd1 vccd1 vccd1 hold1967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1978 _07771_/X vssd1 vssd1 vccd1 vccd1 _14387_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09243__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1989 _14526_/Q vssd1 vssd1 vccd1 vccd1 hold1989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07787_ hold409/X _13725_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold410/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout643_A _15199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09526_ _10166_/A _10338_/B _09979_/C _09979_/D vssd1 vssd1 vccd1 vccd1 _09527_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_91_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08122__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09457_/A _09587_/A _09557_/A _09457_/D vssd1 vssd1 vccd1 vccd1 _09599_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_0_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout810_A _14489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11712__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _09387_/B _09387_/C _09387_/A vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08339_ _08172_/A _08338_/C _08172_/B _08338_/X _07313_/X vssd1 vssd1 vccd1 vccd1
+ _08528_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09622__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11350_ _11351_/B _11620_/B _15221_/Q _11541_/A vssd1 vssd1 vccd1 vccd1 _11352_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11281_ _11281_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11282_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08189__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07637__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ _13020_/A _13020_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _13020_/X sky130_fd_sc_hd__or3b_1
X_10232_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10233_/C sky130_fd_sc_hd__nor2_1
XANTENNA__09925__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__B1 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _10164_/A _10336_/A _10164_/C vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__nor3_1
XANTENNA__10091__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _10246_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10094_/Y sky130_fd_sc_hd__nor2_1
X_14971_ _14971_/CLK _14971_/D vssd1 vssd1 vccd1 vccd1 _14971_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09233__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13922_ _15289_/CLK _13922_/D vssd1 vssd1 vccd1 vccd1 _13922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09153__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13853_ _14612_/CLK hold686/X vssd1 vssd1 vccd1 vccd1 hold685/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ _13393_/B _13104_/A2 _12803_/X vssd1 vssd1 vccd1 vccd1 _12804_/X sky130_fd_sc_hd__a21o_1
X_10996_ _10996_/A _10996_/B _10996_/C _10996_/D vssd1 vssd1 vccd1 vccd1 _10996_/Y
+ sky130_fd_sc_hd__nand4_4
X_13784_ hold259/X vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _14670_/Q _13943_/Q _12735_/S vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__mux2_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13403__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _14344_/Q _14248_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _12666_/X sky130_fd_sc_hd__mux2_1
X_15454_ _15454_/CLK hold716/X vssd1 vssd1 vccd1 vccd1 hold715/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13096__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11617_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14405_ _15438_/CLK hold782/X vssd1 vssd1 vccd1 vccd1 hold781/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ _14792_/Q _14504_/Q _14632_/Q _14728_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12597_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_68_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15385_ _15385_/CLK _15385_/D vssd1 vssd1 vccd1 vccd1 _15385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10759__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ _11548_/A _11548_/B vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__xnor2_1
X_14336_ _14750_/CLK hold338/X vssd1 vssd1 vccd1 vccd1 hold337/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold508 hold508/A vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold519 hold519/A vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ _15360_/CLK hold510/X vssd1 vssd1 vccd1 vccd1 hold509/A sky130_fd_sc_hd__dfxtp_1
X_11479_ _11479_/A _11479_/B vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ hold927/X _13664_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 hold928/A sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11577__B _14970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14198_ _15087_/CLK _14198_/D vssd1 vssd1 vccd1 vccd1 _14198_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08275__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13389_/A _13149_/B vssd1 vssd1 vccd1 vccd1 _15014_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 _06988_/X vssd1 vssd1 vccd1 vccd1 _13807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1219 _14329_/Q vssd1 vssd1 vccd1 vccd1 hold1219/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09224__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08886__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ _13683_/A _11729_/B _07744_/A vssd1 vssd1 vccd1 vccd1 _07710_/X sky130_fd_sc_hd__and3b_4
XFILLER_0_75_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08690_ _08689_/A _08689_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08691_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_205_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07641_ hold1441/X _13714_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_205_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15215__D _15215_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _13396_/A _07572_/B vssd1 vssd1 vccd1 vccd1 _14197_/D sky130_fd_sc_hd__and2_1
XANTENNA__12436__B1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08104__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ _09178_/Y _09180_/X _09309_/Y _09310_/X vssd1 vssd1 vccd1 vccd1 _09314_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_165_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12987__A1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10937__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09242_ _09227_/Y _09232_/Y _09241_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09243_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10656__B _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07311__A _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _09173_/A _09297_/B _09173_/C vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_173_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ hold337/A hold913/A _14400_/Q _14112_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _08125_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11411__A1 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11411__B2 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ hold893/A _15266_/Q _15074_/Q _14367_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08055_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07006_ _13744_/A1 hold2235/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07006_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09238__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12598__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__A _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2410 _14831_/Q vssd1 vssd1 vccd1 vccd1 hold2410/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput106 in1[18] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput117 in1[28] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_1
Xhold2421 _12093_/X vssd1 vssd1 vccd1 vccd1 _14858_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07981__A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput128 in1[9] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_1
Xhold2432 _14051_/Q vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xinput139 in2[19] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _09119_/A _08957_/B vssd1 vssd1 vccd1 vccd1 _08957_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout760_A _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2443 _13467_/X vssd1 vssd1 vccd1 vccd1 _15227_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2454 hold2852/X vssd1 vssd1 vccd1 vccd1 _06903_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13467__A2 _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout858_A _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1720 _13704_/X vssd1 vssd1 vccd1 vccd1 _15410_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11707__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2465 _14867_/Q vssd1 vssd1 vccd1 vccd1 hold2465/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2476 _12107_/X vssd1 vssd1 vccd1 vccd1 _14865_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07908_ _07908_/A _07908_/B _07908_/C vssd1 vssd1 vccd1 vccd1 _07908_/X sky130_fd_sc_hd__and3_1
Xhold1731 _15284_/Q vssd1 vssd1 vccd1 vccd1 hold1731/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _09253_/A _09435_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _08888_/X sky130_fd_sc_hd__and3_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2487 _14845_/Q vssd1 vssd1 vccd1 vccd1 hold2487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1742 _07145_/X vssd1 vssd1 vccd1 vccd1 _13955_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2498 _15347_/Q vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__clkbuf_2
Xhold1753 _14495_/Q vssd1 vssd1 vccd1 vccd1 hold1753/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1764 _11673_/X vssd1 vssd1 vccd1 vccd1 _14476_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07192__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1775 _13979_/Q vssd1 vssd1 vccd1 vccd1 hold1775/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _07862_/C _14031_/Q _14034_/Q _06909_/Y vssd1 vssd1 vccd1 vccd1 _07839_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_196_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1786 _11739_/X vssd1 vssd1 vccd1 vccd1 _14533_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1797 _14782_/Q vssd1 vssd1 vccd1 vccd1 hold1797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _10850_/A _10850_/B _10850_/C vssd1 vssd1 vccd1 vccd1 _10850_/X sky130_fd_sc_hd__and3_2
XFILLER_0_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13624__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _14349_/Q _14253_/Q hold475/A _14125_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09510_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12978__B2 _13198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10781_ _14967_/Q _10781_/B vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__and2_1
XFILLER_0_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _12520_/A _12520_/B _12601_/A vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__or3b_1
XANTENNA__10453__A2 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08317__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12676_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12452_/C sky130_fd_sc_hd__or2_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12825__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15170_ _15268_/CLK _15170_/D vssd1 vssd1 vccd1 vccd1 _15170_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12382_ _07919_/B _08636_/Y _13142_/B _13081_/A1 _13455_/A vssd1 vssd1 vccd1 vccd1
+ _14943_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_90 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _14409_/CLK hold858/X vssd1 vssd1 vccd1 vccd1 hold857/A sky130_fd_sc_hd__dfxtp_1
X_11333_ _11526_/A _11333_/B _15223_/Q _15224_/Q vssd1 vssd1 vccd1 vccd1 _11334_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _15422_/CLK _14052_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12589__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ _11460_/A _11264_/B _11328_/B _11264_/D vssd1 vssd1 vccd1 vccd1 _11460_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13003_ _13711_/A1 _13103_/A2 _13078_/B1 _13199_/B vssd1 vssd1 vccd1 vccd1 _13003_/X
+ sky130_fd_sc_hd__a22o_1
X_10215_ _10392_/A _10213_/X _09970_/Y _09973_/Y vssd1 vssd1 vccd1 vccd1 _10215_/X
+ sky130_fd_sc_hd__o211a_1
X_11195_ _11564_/A _11378_/D _11196_/C _11382_/A vssd1 vssd1 vccd1 vccd1 _11195_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08987__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _10007_/X _10011_/B _10312_/B _10145_/X vssd1 vssd1 vccd1 vccd1 _10148_/B
+ sky130_fd_sc_hd__o211ai_2
X_10077_ _12221_/B _10077_/B vssd1 vssd1 vccd1 vccd1 _10077_/Y sky130_fd_sc_hd__nand2_1
X_14954_ _14954_/CLK _14954_/D vssd1 vssd1 vccd1 vccd1 _14954_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _15438_/CLK _13905_/D vssd1 vssd1 vccd1 vccd1 _13905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ _14989_/CLK _14885_/D vssd1 vssd1 vccd1 vccd1 _14885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08885__A2 _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09509__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ _14595_/CLK _13836_/D vssd1 vssd1 vccd1 vccd1 _13836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11316__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12969__A1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10979_ _11569_/A _11606_/B _11570_/B _11563_/A vssd1 vssd1 vccd1 vccd1 _10979_/X
+ sky130_fd_sc_hd__a22o_1
X_13767_ hold253/X vssd1 vssd1 vccd1 vccd1 hold254/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12718_ _12749_/S1 _12715_/X _12717_/X vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10476__B _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13698_ hold909/X _13698_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 hold910/A sky130_fd_sc_hd__mux2_1
XFILLER_0_128_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15437_ _15437_/CLK hold766/X vssd1 vssd1 vccd1 vccd1 hold765/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ _13875_/Q _14003_/Q _13843_/Q _13811_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12649_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _15416_/CLK _15368_/D vssd1 vssd1 vccd1 vccd1 _15368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11588__A _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14319_ _15379_/CLK _14319_/D vssd1 vssd1 vccd1 vccd1 _14319_/Q sky130_fd_sc_hd__dfxtp_1
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15299_ _15299_/CLK _15299_/D vssd1 vssd1 vccd1 vccd1 _15299_/Q sky130_fd_sc_hd__dfxtp_1
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold338 hold338/A vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 hold349/A vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09860_ _09860_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__nand2_2
XANTENNA__10642__D _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout807 _12365_/S1 vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout818 _14489_/Q vssd1 vssd1 vccd1 vccd1 _13098_/S1 sky130_fd_sc_hd__buf_4
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 _14488_/Q vssd1 vssd1 vccd1 vccd1 _12365_/S0 sky130_fd_sc_hd__buf_4
XANTENNA__08573__A1 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _08926_/A _09864_/A _08810_/C _08922_/A vssd1 vssd1 vccd1 vccd1 _08812_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08573__B2 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _14802_/Q _14514_/Q hold323/A hold865/A _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09792_/B sky130_fd_sc_hd__mux4_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _14750_/Q vssd1 vssd1 vccd1 vccd1 hold1005/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 _11877_/X vssd1 vssd1 vccd1 vccd1 _14699_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13308__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1027 _14109_/Q vssd1 vssd1 vccd1 vccd1 hold1027/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _09346_/B _08743_/C _08743_/A vssd1 vssd1 vccd1 vccd1 _08742_/X sky130_fd_sc_hd__o21a_1
Xhold1038 _11890_/X vssd1 vssd1 vccd1 vccd1 _14712_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _14212_/Q vssd1 vssd1 vccd1 vccd1 hold1049/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12212__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__A _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08673_ _08673_/A _08673_/B vssd1 vssd1 vccd1 vccd1 _08674_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_206_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_186_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15264_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13742__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ hold1835/X _13730_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07624_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_178_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07740__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07555_ _13393_/A _07555_/B vssd1 vssd1 vccd1 vccd1 _14180_/D sky130_fd_sc_hd__and2_1
XANTENNA__09825__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09825__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _07512_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ hold2814/X hold285/X _07493_/S vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__mux2_1
XFILLER_0_36_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09225_ _13879_/Q hold291/A _13847_/Q _13815_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09225_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout606_A _15209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _09027_/A _09027_/B _09027_/C vssd1 vssd1 vccd1 vccd1 _09157_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08107_ _08107_/A hold443/X vssd1 vssd1 vccd1 vccd1 _08108_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _09087_/A _09087_/B _09087_/C vssd1 vssd1 vccd1 vccd1 _09350_/C sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_110_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15090_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07187__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ _08038_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08039_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold850 hold850/A vssd1 vssd1 vccd1 vccd1 hold850/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12106__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 hold861/A vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__C1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__B _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 hold872/A vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 hold883/A vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 hold894/A vssd1 vssd1 vccd1 vccd1 hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _10000_/A _11578_/A _10108_/C _14963_/Q vssd1 vssd1 vccd1 vccd1 _10000_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__08564__A1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07998__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _09831_/B _09833_/B _09986_/X _09988_/Y vssd1 vssd1 vccd1 vccd1 _09989_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2240 _11736_/X vssd1 vssd1 vccd1 vccd1 _14530_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2251 _14458_/Q vssd1 vssd1 vccd1 vccd1 hold2251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2262 _13506_/X vssd1 vssd1 vccd1 vccd1 _15264_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12122__A _15001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2273 _13905_/Q vssd1 vssd1 vccd1 vccd1 hold2273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08316__A1 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2284 _13477_/X vssd1 vssd1 vccd1 vccd1 _15236_/D sky130_fd_sc_hd__buf_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2295 _15274_/Q vssd1 vssd1 vccd1 vccd1 hold2295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 _07097_/X vssd1 vssd1 vccd1 vccd1 _13910_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1561 _14354_/Q vssd1 vssd1 vccd1 vccd1 hold1561/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_177_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15438_/CLK sky130_fd_sc_hd__clkbuf_16
X_11951_ _13739_/A1 hold1363/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11951_/X sky130_fd_sc_hd__mux2_1
Xhold1572 _07142_/X vssd1 vssd1 vccd1 vccd1 _13952_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1583 _14791_/Q vssd1 vssd1 vccd1 vccd1 hold1583/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1594 _07759_/X vssd1 vssd1 vccd1 vccd1 _14375_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13652__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _10675_/Y _10719_/X _11085_/B _10901_/Y vssd1 vssd1 vccd1 vccd1 _11091_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14670_ _15056_/CLK _14670_/D vssd1 vssd1 vccd1 vccd1 _14670_/Q sky130_fd_sc_hd__dfxtp_1
X_11882_ hold1041/X _13703_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 _11882_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07650__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13621_ input36/X _13636_/B vssd1 vssd1 vccd1 vccd1 _13621_/X sky130_fd_sc_hd__or2_1
X_10833_ _10830_/Y _10831_/X _10642_/X _10645_/X vssd1 vssd1 vccd1 vccd1 _10834_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__B _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13552_ _14432_/Q _13554_/B vssd1 vssd1 vccd1 vccd1 _13552_/X sky130_fd_sc_hd__or2_1
X_10764_ _11504_/A _10761_/X _10763_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _10765_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _13724_/A1 _12329_/B _12953_/B1 _13179_/B vssd1 vssd1 vccd1 vccd1 _12503_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13483_ _13487_/A hold107/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__and2_1
XFILLER_0_192_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ _10482_/A _10481_/B _10479_/X vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11900__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15222_ _15222_/CLK _15222_/D vssd1 vssd1 vccd1 vccd1 _15222_/Q sky130_fd_sc_hd__dfxtp_4
X_12434_ hold661/X hold2209/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12434_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09044__A2 _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15153_ _15316_/CLK _15153_/D vssd1 vssd1 vccd1 vccd1 _15153_/Q sky130_fd_sc_hd__dfxtp_1
X_12365_ hold275/A hold301/A _14591_/Q _13960_/Q _12365_/S0 _12365_/S1 vssd1 vssd1
+ vccd1 vccd1 _12366_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_121_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_101_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15244_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07097__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14104_ _14105_/CLK hold268/X vssd1 vssd1 vccd1 vccd1 _14104_/Q sky130_fd_sc_hd__dfxtp_1
X_11316_ hold783/A _14555_/Q hold655/A hold795/A _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _11316_/X sky130_fd_sc_hd__mux4_1
X_15084_ _15373_/CLK _15084_/D vssd1 vssd1 vccd1 vccd1 _15084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12296_ _07439_/A _14088_/Q _11729_/C _15350_/Q _12295_/X vssd1 vssd1 vccd1 vccd1
+ _12296_/X sky130_fd_sc_hd__a221o_1
XANTENNA_output260_A _14877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ _15425_/CLK _14035_/D vssd1 vssd1 vccd1 vccd1 _14035_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _11517_/A _15221_/Q _11247_/C _11348_/A vssd1 vssd1 vccd1 vccd1 _11348_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08004__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11177_/B _11177_/C _11177_/A vssd1 vssd1 vccd1 vccd1 _11179_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10129_ _10129_/A _10827_/D vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13300__A1 input139/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12103__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ _15389_/CLK _14937_/D vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_168_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15373_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08858__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14868_ _14876_/CLK _14868_/D vssd1 vssd1 vccd1 vccd1 _14868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__C _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11590__B _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13819_ _15378_/CLK _13819_/D vssd1 vssd1 vccd1 vccd1 _13819_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10487__A _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14799_ _15376_/CLK _14799_/D vssd1 vssd1 vccd1 vccd1 _14799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07340_ _07849_/B vssd1 vssd1 vccd1 vccd1 _07341_/B sky130_fd_sc_hd__inv_2
XFILLER_0_35_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12811__B1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A2 _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07271_ _07271_/A _09340_/A vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10637__D _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ _09253_/A _09712_/B _09011_/C _09011_/D vssd1 vssd1 vccd1 vccd1 _09010_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__11810__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2738_A _15182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13737__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _09912_/A _11283_/S vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__or2_1
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12641__S _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout604 _15209_/Q vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12878__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout615 _15206_/Q vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__buf_6
XFILLER_0_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout626 _10033_/A vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07735__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12973__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _09690_/B _09692_/B _09841_/X _09842_/Y vssd1 vssd1 vccd1 vccd1 _09896_/A
+ sky130_fd_sc_hd__a211oi_4
Xfanout637 _08012_/B vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__buf_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout648 _15198_/Q vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__buf_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout659 hold2794/X vssd1 vssd1 vccd1 vccd1 _13746_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout389_A _11652_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _13691_/A1 hold745/X _06994_/S vssd1 vssd1 vccd1 vccd1 hold746/A sky130_fd_sc_hd__mux2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__nand2_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12725__S0 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ _08725_/A _08725_/B _08621_/B vssd1 vssd1 vccd1 vccd1 _08725_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_159_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _14569_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_174_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12877__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout556_A _15423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08760_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _08656_/Y sky130_fd_sc_hd__nor2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08793__C _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07607_ _13746_/A1 hold2113/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07607_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08586_/B _08586_/C _08586_/A vssd1 vssd1 vccd1 vccd1 _08589_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10397__A _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout723_A _14962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ hold477/X _13742_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold478/A sky130_fd_sc_hd__mux2_1
XFILLER_0_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ hold145/X _07475_/B vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__and2_1
XFILLER_0_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11720__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ _11473_/A _09203_/Y _09204_/X _09207_/X vssd1 vssd1 vccd1 vccd1 _13390_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__13501__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10480_ _10477_/Y _10478_/X _10303_/X _10305_/X vssd1 vssd1 vccd1 vccd1 _10481_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_112_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _09138_/A _09866_/B _09138_/C _09138_/D vssd1 vssd1 vccd1 vccd1 _09139_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12150_ _14886_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__D _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _10959_/X _10960_/X _11099_/Y _11281_/B _10397_/A vssd1 vssd1 vccd1 vccd1
+ _11101_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ hold2448/X _12099_/A2 _12080_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12081_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10860__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_127_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 hold680/A vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold691 hold691/A vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07645__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11032_ _11029_/X _11030_/Y _10847_/X _10850_/X vssd1 vssd1 vccd1 vccd1 _11033_/D
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09426__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12964__S0 _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2070 _07592_/X vssd1 vssd1 vccd1 vccd1 _14216_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2081 _13908_/Q vssd1 vssd1 vccd1 vccd1 hold2081/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2092 _07064_/X vssd1 vssd1 vccd1 vccd1 _13880_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ hold1659/X hold869/X hold1037/X hold773/X _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12983_/X sky130_fd_sc_hd__mux4_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1380 _11863_/X vssd1 vssd1 vccd1 vccd1 _14685_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _15042_/CLK _14722_/D vssd1 vssd1 vccd1 vccd1 _14722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1391 _14243_/Q vssd1 vssd1 vccd1 vccd1 hold1391/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10647__A2 _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ _13689_/A1 hold1167/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _15427_/CLK _14653_/D vssd1 vssd1 vccd1 vccd1 _14653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ hold1253/X _13719_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ input58/X _13625_/B _13625_/C vssd1 vssd1 vccd1 vccd1 _15329_/D sky130_fd_sc_hd__and3_1
XFILLER_0_184_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10816_ _10817_/A _10817_/B _10817_/C vssd1 vssd1 vccd1 vccd1 _10816_/X sky130_fd_sc_hd__and3_1
XANTENNA__10100__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14584_ _14926_/CLK hold158/X vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
X_11796_ _13716_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__09265__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13535_ _13535_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _15293_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _10568_/B _10405_/B _10744_/A vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13411__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ _11526_/A _11550_/A _15219_/Q _11620_/B vssd1 vssd1 vccd1 vccd1 _10681_/A
+ sky130_fd_sc_hd__nand4_1
X_13466_ _13466_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _13466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09648__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15205_ _15324_/CLK _15205_/D vssd1 vssd1 vccd1 vccd1 _15205_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_106_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12417_ _12642_/A1 _12416_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12417_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12027__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ _13397_/A _13397_/B vssd1 vssd1 vccd1 vccd1 _15188_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10473__C _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10032__B1 _14957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput207 _14171_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[1] sky130_fd_sc_hd__buf_12
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput218 _14172_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[2] sky130_fd_sc_hd__buf_12
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15136_ _15304_/CLK _15136_/D vssd1 vssd1 vccd1 vccd1 _15136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput229 _14434_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[10] sky130_fd_sc_hd__buf_12
X_12348_ _14622_/Q _14718_/Q _12466_/S vssd1 vssd1 vccd1 vccd1 _12348_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12279_ _13168_/A _13444_/B vssd1 vssd1 vccd1 vccd1 _14928_/D sky130_fd_sc_hd__nor2_2
X_15067_ _15384_/CLK _15067_/D vssd1 vssd1 vccd1 vccd1 _15067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _14483_/CLK hold294/X vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08510_ _08511_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08510_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11805__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10638__A2 _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09490_ _09491_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__nand2b_1
XProc_895 vssd1 vssd1 vccd1 vccd1 imemreq_val Proc_895/LO sky130_fd_sc_hd__conb_1
XFILLER_0_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__A1 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08441_ _13554_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08441_/X sky130_fd_sc_hd__or2_1
XANTENNA_hold2590_A _12270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07303__B _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ _06926_/A _08365_/Y _08367_/Y _08369_/Y _08371_/Y vssd1 vssd1 vccd1 vccd1
+ _08372_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07323_ _07323_/A _07323_/B _07323_/C _07887_/A vssd1 vssd1 vccd1 vccd1 _07330_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _15224_/Q _14968_/Q vssd1 vssd1 vccd1 vccd1 _07255_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10249__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ hold1101/X _13653_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07185_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_171_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10574__A1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07973__B _07974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10680__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _07477_/Y vssd1 vssd1 vccd1 vccd1 _07493_/S sky130_fd_sc_hd__buf_12
XANTENNA__09246__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12946__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 _07080_/Y vssd1 vssd1 vccd1 vccd1 _07112_/S sky130_fd_sc_hd__buf_8
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout423 _11961_/Y vssd1 vssd1 vccd1 vccd1 _11977_/S sky130_fd_sc_hd__clkbuf_16
Xfanout434 _07778_/Y vssd1 vssd1 vccd1 vccd1 _07810_/S sky130_fd_sc_hd__clkbuf_16
Xfanout445 _07389_/Y vssd1 vssd1 vccd1 vccd1 _13797_/A2 sky130_fd_sc_hd__buf_4
Xfanout456 _07012_/Y vssd1 vssd1 vccd1 vccd1 _07044_/S sky130_fd_sc_hd__clkbuf_16
X_09826_ _10183_/A _09979_/B _11588_/A _11623_/A vssd1 vssd1 vccd1 vccd1 _09828_/D
+ sky130_fd_sc_hd__nand4_1
Xfanout467 _11287_/S vssd1 vssd1 vccd1 vccd1 _12221_/B sky130_fd_sc_hd__buf_8
Xfanout478 _07355_/Y vssd1 vssd1 vccd1 vccd1 _13081_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout489 _12126_/B vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09757_ _09754_/X _09755_/Y _09608_/X _09610_/Y vssd1 vssd1 vccd1 vccd1 _09758_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout840_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06969_ _14084_/Q _14085_/Q _14091_/Q vssd1 vssd1 vccd1 vccd1 _06970_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11715__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _08805_/A _08707_/C _08707_/A vssd1 vssd1 vccd1 vccd1 _08709_/C sky130_fd_sc_hd__a21o_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11826__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09549_/X _09551_/Y _09686_/X _09687_/Y vssd1 vssd1 vccd1 vccd1 _09690_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08640_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08639_/X sky130_fd_sc_hd__and2_1
XANTENNA__13028__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ _13598_/A _11650_/B vssd1 vssd1 vccd1 vccd1 _11650_/Y sky130_fd_sc_hd__nor2_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09247__A2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _10601_/A _10952_/A vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__or2_1
XFILLER_0_182_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _11581_/A _11581_/B vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12251__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13320_ _13338_/A _13320_/B vssd1 vssd1 vccd1 vccd1 _15126_/D sky130_fd_sc_hd__nor2_1
X_10532_ _10532_/A _10532_/B _10532_/C vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13251_ _13287_/A _13251_/B vssd1 vssd1 vccd1 vccd1 _15103_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_190_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10463_ _10463_/A _10463_/B _10463_/C vssd1 vssd1 vccd1 vccd1 _10464_/C sky130_fd_sc_hd__nor3_1
XFILLER_0_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11389__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12554__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ hold589/A hold289/A hold855/A _14717_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12202_/X sky130_fd_sc_hd__mux4_1
X_13182_ _13481_/A _13182_/B vssd1 vssd1 vccd1 vccd1 _15047_/D sky130_fd_sc_hd__and2_1
X_10394_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10565__A1 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__A0 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12133_ _12066_/A _12195_/A2 _12132_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09707__B1 _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _14097_/Q _14096_/Q _14095_/Q vssd1 vssd1 vccd1 vccd1 _12124_/D sky130_fd_sc_hd__or3b_2
XANTENNA__10317__A1 _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11514__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _11015_/A _11015_/B vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__or2_1
XFILLER_0_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08210__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13406__A _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _14356_/Q hold433/X _13066_/S vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _15410_/CLK hold934/X vssd1 vssd1 vccd1 vccd1 hold933/A sky130_fd_sc_hd__dfxtp_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _15058_/Q hold865/X _11927_/S vssd1 vssd1 vccd1 vccd1 hold866/A sky130_fd_sc_hd__mux2_1
XFILLER_0_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _14804_/Q hold649/A hold847/A _14740_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12897_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08219__B _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10468__C _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _15179_/CLK _14636_/D vssd1 vssd1 vccd1 vccd1 _14636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11848_ hold1335/X _13735_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 _11848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10765__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ _15079_/CLK hold230/X vssd1 vssd1 vccd1 vccd1 hold229/A sky130_fd_sc_hd__dfxtp_1
X_11779_ hold1437/X _13666_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13141__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13518_ _13666_/A1 hold947/X _13518_/S vssd1 vssd1 vccd1 vccd1 hold948/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ _15042_/CLK hold790/X vssd1 vssd1 vccd1 vccd1 hold789/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13449_ _09919_/B _13450_/A _13448_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15218_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08749__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13742__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11596__A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15119_ _15127_/CLK _15119_/D vssd1 vssd1 vccd1 vccd1 _15119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08990_ hold609/A _14540_/Q hold737/A _14764_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08990_/X sky130_fd_sc_hd__mux4_1
Xhold2806 _12739_/X vssd1 vssd1 vccd1 vccd1 hold2806/X sky130_fd_sc_hd__dlygate4sd3_1
X_07941_ hold957/A _13929_/Q _15430_/Q _13897_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07942_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2817 _15067_/Q vssd1 vssd1 vccd1 vccd1 hold2817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2828 _15320_/Q vssd1 vssd1 vccd1 vccd1 hold2828/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15218__D _15218_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2839 _15300_/Q vssd1 vssd1 vccd1 vccd1 hold2839/X sky130_fd_sc_hd__dlygate4sd3_1
X_07872_ _07862_/A _14088_/Q _11729_/C _15345_/Q _07871_/X vssd1 vssd1 vccd1 vccd1
+ _07872_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_103_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09611_ _09608_/X _09609_/Y _09394_/X _09397_/X vssd1 vssd1 vccd1 vccd1 _09611_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09542_ _09542_/A _09979_/B _15209_/Q _09860_/B vssd1 vssd1 vccd1 vccd1 _09673_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__07314__A _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09473_ _09328_/Y _09330_/Y _09471_/X _09472_/Y vssd1 vssd1 vccd1 vccd1 _09760_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12481__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15256_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ _08329_/A _08329_/C _08329_/B vssd1 vssd1 vccd1 vccd1 _08427_/C sky130_fd_sc_hd__a21boi_1
XFILLER_0_164_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12769__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08355_ hold225/A _14307_/Q _14598_/Q _13967_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08355_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_4_9__f_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout421_A _13204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07306_ _08702_/B _11541_/A vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout519_A _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13051__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08286_ hold2750/X input31/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13180_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07237_ _07237_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07660__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09937__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ _13669_/A1 hold1847/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout790_A _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A2 _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout888_A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07099_ _13735_/A1 hold1667/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07099_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07195__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12114__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08373__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09809_ _10166_/A _10338_/B _09809_/C _11536_/B vssd1 vssd1 vccd1 vccd1 _09964_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_92_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ _12820_/A _12820_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12827_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_201_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12951_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _12752_/C sky130_fd_sc_hd__or2_1
XFILLER_0_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13660__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15454_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ hold789/X _13656_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold790/A sky130_fd_sc_hd__mux2_1
XFILLER_0_167_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _13150_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _14955_/D sky130_fd_sc_hd__nor2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14776_/CLK hold310/X vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__dfxtp_1
X_11633_ _11633_/A _11633_/B vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12224__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10585__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14352_ _15196_/CLK hold932/X vssd1 vssd1 vccd1 vccd1 hold931/A sky130_fd_sc_hd__dfxtp_1
X_11564_ _11564_/A _11564_/B vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ input141/X fanout5/X fanout3/X input109/X vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__a22o_1
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__or2_1
XFILLER_0_135_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11495_ _11497_/A _11495_/B vssd1 vssd1 vccd1 vccd1 _11495_/Y sky130_fd_sc_hd__nor2_1
X_14283_ _15444_/CLK _14283_/D vssd1 vssd1 vccd1 vccd1 _14283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09928__B1 _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10446_ _10629_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10464_/A sky130_fd_sc_hd__or2_1
X_13234_ hold753/X _13680_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold754/A sky130_fd_sc_hd__mux2_1
XANTENNA_output173_A _15166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ _10196_/Y _10199_/Y _10439_/A _10376_/X vssd1 vssd1 vccd1 vccd1 _10439_/B
+ sky130_fd_sc_hd__a211oi_2
X_13165_ _13390_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _15030_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _14998_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12116_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_23_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13096_ hold367/A hold769/A hold535/A _14393_/Q _13091_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13096_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12047_ _12059_/A _12047_/B vssd1 vssd1 vccd1 vccd1 _14836_/D sky130_fd_sc_hd__and2_1
XFILLER_0_100_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13136__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _14783_/CLK hold422/X vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__dfxtp_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12463__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _13887_/Q _14015_/Q hold739/A hold761/A _12915_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12949_/X sky130_fd_sc_hd__mux4_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15068_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_191 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14619_ _15063_/CLK hold354/X vssd1 vssd1 vccd1 vccd1 hold353/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _08312_/A _09138_/A vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10777__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08071_ hold2729/X input28/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13177_/B sky130_fd_sc_hd__mux2_2
XANTENNA_hold2553_A _14995_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ hold1701/X _13512_/A0 _07028_/S vssd1 vssd1 vccd1 vccd1 _07022_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13715__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10529__A1 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10434__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07954__D _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2603 _12149_/X vssd1 vssd1 vccd1 vccd1 _14885_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08973_ _09087_/B _09222_/B vssd1 vssd1 vccd1 vccd1 _08973_/X sky130_fd_sc_hd__or2_1
Xhold2614 hold2828/X vssd1 vssd1 vccd1 vccd1 _10744_/B sky130_fd_sc_hd__clkbuf_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2625 _14888_/Q vssd1 vssd1 vccd1 vccd1 _12154_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13745__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2636 _15329_/Q vssd1 vssd1 vccd1 vccd1 _07345_/A sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _14426_/Q _13591_/A2 _07926_/A _07923_/Y vssd1 vssd1 vccd1 vccd1 _07924_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2647 hold2831/X vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__clkbuf_2
Xhold1902 _07159_/X vssd1 vssd1 vccd1 vccd1 _13967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2658 _14821_/Q vssd1 vssd1 vccd1 vccd1 hold2658/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12845__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1913 _13891_/Q vssd1 vssd1 vccd1 vccd1 hold1913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1924 _11747_/X vssd1 vssd1 vccd1 vccd1 _14541_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2669 _12006_/X vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09524__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1935 _13806_/Q vssd1 vssd1 vccd1 vccd1 hold1935/X sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _07855_/A _07857_/C _07855_/C vssd1 vssd1 vccd1 vccd1 _11283_/S sky130_fd_sc_hd__or3_4
XFILLER_0_78_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1946 _11964_/X vssd1 vssd1 vccd1 vccd1 _14783_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10701__A1 _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1957 _13954_/Q vssd1 vssd1 vccd1 vccd1 hold1957/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1968 _07773_/X vssd1 vssd1 vccd1 vccd1 _14389_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout469_A _07884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1979 _13935_/Q vssd1 vssd1 vccd1 vccd1 hold1979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07786_ hold441/X _13724_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold442/A sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09525_ _10338_/B _09979_/C _09979_/D _10166_/A vssd1 vssd1 vccd1 vccd1 _09527_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12454__A1 _13379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12995__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14876_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08753__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09453_/Y _09454_/X _09270_/Y _09273_/X vssd1 vssd1 vccd1 vccd1 _09457_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08598_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_149_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12206__A1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09387_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout803_A _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ _08702_/B _11541_/A _08338_/C vssd1 vssd1 vccd1 vccd1 _08338_/X sky130_fd_sc_hd__and3_1
XFILLER_0_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__A2 _13393_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08269_ _08873_/A _08266_/X _08268_/X vssd1 vssd1 vccd1 vccd1 _08269_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10300_ _11620_/A _11537_/B vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ _11280_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08603__A _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__and2_1
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11193__A1 _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__B2 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _10336_/A _10164_/C _10164_/A vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_207_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13655__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14970_ _15418_/CLK _14970_/D vssd1 vssd1 vccd1 vccd1 _14970_/Q sky130_fd_sc_hd__dfxtp_2
X_10093_ _10426_/A _10090_/X _10092_/X _10255_/A1 vssd1 vssd1 vccd1 vccd1 _10094_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09233__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07653__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13921_ _15454_/CLK _13921_/D vssd1 vssd1 vccd1 vccd1 _13921_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12693__A1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09153__B _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ _15191_/CLK _13852_/D vssd1 vssd1 vccd1 vccd1 _13852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12803_ _13736_/A1 _13103_/A2 _13078_/B1 _13191_/B vssd1 vssd1 vccd1 vccd1 _12803_/X
+ sky130_fd_sc_hd__a22o_1
X_13783_ hold157/X vssd1 vssd1 vccd1 vccd1 hold158/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15356_/CLK sky130_fd_sc_hd__clkbuf_16
X_10995_ _10994_/B _10994_/C _10994_/A vssd1 vssd1 vccd1 vccd1 _10996_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11903__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08113__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07889__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12734_ hold723/A _13911_/Q _12735_/S vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__mux2_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15453_/CLK hold834/X vssd1 vssd1 vccd1 vccd1 hold833/A sky130_fd_sc_hd__dfxtp_1
X_12665_ hold1833/X hold1811/X _12665_/S vssd1 vssd1 vccd1 vccd1 _12665_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07872__B2 _15345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14404_ _14955_/CLK hold960/X vssd1 vssd1 vccd1 vccd1 hold959/A sky130_fd_sc_hd__dfxtp_1
X_11616_ _11626_/B _11397_/B _11397_/C _11401_/A vssd1 vssd1 vccd1 vccd1 _11617_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15384_ _15384_/CLK hold316/X vssd1 vssd1 vccd1 vccd1 hold315/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12596_ hold471/A hold705/A hold981/A _14373_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12596_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11956__A0 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10759__A1 _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14335_ _15391_/CLK hold416/X vssd1 vssd1 vccd1 vccd1 hold415/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11547_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11548_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12734__S _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 hold509/A vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14266_ _15263_/CLK hold620/X vssd1 vssd1 vccd1 vccd1 hold619/A sky130_fd_sc_hd__dfxtp_1
X_11478_ _11645_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11479_/B sky130_fd_sc_hd__or2_1
XFILLER_0_204_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13217_ hold2097/X _13663_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__mux2_1
X_10429_ hold419/A hold983/A hold331/A _14774_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10429_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14197_ _15190_/CLK _14197_/D vssd1 vssd1 vccd1 vccd1 _14197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13150_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _15013_/D sky130_fd_sc_hd__nor2_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__A1 _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _11474_/X _13104_/A2 _13078_/X vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1209 _14365_/Q vssd1 vssd1 vccd1 vccd1 hold1209/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09224__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07640_ hold797/X _13680_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold798/A sky130_fd_sc_hd__mux2_1
XFILLER_0_205_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07571_ _13396_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _14196_/D sky130_fd_sc_hd__and2_1
XANTENNA__12436__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12909__S _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15199_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08104__A2 _13379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ _09307_/X _09308_/Y _09175_/B _09178_/B vssd1 vssd1 vccd1 vccd1 _09310_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11813__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09241_ _10430_/B1 _09234_/Y _09236_/Y _09238_/Y _09240_/Y vssd1 vssd1 vccd1 vccd1
+ _09241_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_111_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2768_A _15194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15231__D _15231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ _10185_/A _09858_/C _09171_/C _09297_/A vssd1 vssd1 vccd1 vccd1 _09173_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07311__B _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11947__A0 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08123_ _08760_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _08123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_146_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11411__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08197_/A _08051_/X _08053_/X vssd1 vssd1 vccd1 vccd1 _08054_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07738__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09519__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07005_ hold2765/A hold2193/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07005_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12598__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08142__B _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2400 _15307_/Q vssd1 vssd1 vccd1 vccd1 _08851_/A sky130_fd_sc_hd__buf_1
Xinput107 in1[19] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_1
Xhold2411 _12036_/X vssd1 vssd1 vccd1 vccd1 _12037_/B sky130_fd_sc_hd__dlygate4sd3_1
Xinput118 in1[29] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__clkbuf_1
Xhold2422 _14857_/Q vssd1 vssd1 vccd1 vccd1 hold2422/X sky130_fd_sc_hd__dlygate4sd3_1
X_08956_ _08840_/A _08842_/B _08840_/B vssd1 vssd1 vccd1 vccd1 _08957_/B sky130_fd_sc_hd__o21ba_1
Xinput129 in2[0] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_2
Xhold2433 _14851_/Q vssd1 vssd1 vccd1 vccd1 hold2433/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2444 hold2854/X vssd1 vssd1 vccd1 vccd1 _10921_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2455 _14866_/Q vssd1 vssd1 vccd1 vccd1 hold2455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1710 _07757_/X vssd1 vssd1 vccd1 vccd1 _14373_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2466 _12111_/X vssd1 vssd1 vccd1 vccd1 _14867_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07907_ _07908_/B _07908_/C vssd1 vssd1 vccd1 vccd1 _07907_/X sky130_fd_sc_hd__and2_1
Xhold1721 _13951_/Q vssd1 vssd1 vccd1 vccd1 hold1721/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1732 _13526_/X vssd1 vssd1 vccd1 vccd1 _15284_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08879__B1 _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2477 _15154_/Q vssd1 vssd1 vccd1 vccd1 hold2477/X sky130_fd_sc_hd__dlygate4sd3_1
X_08887_ _09435_/A _09858_/A _09858_/B _09253_/A vssd1 vssd1 vccd1 vccd1 _08887_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1743 _13917_/Q vssd1 vssd1 vccd1 vccd1 hold1743/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2488 _12067_/X vssd1 vssd1 vccd1 vccd1 _14845_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09540__A1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2499 _14448_/Q vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__buf_1
Xhold1754 _11699_/X vssd1 vssd1 vccd1 vccd1 _14495_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09540__B2 _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1765 _15419_/Q vssd1 vssd1 vccd1 vccd1 hold1765/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ _15343_/Q hold277/A vssd1 vssd1 vccd1 vccd1 _07838_/Y sky130_fd_sc_hd__xnor2_1
Xhold1776 _07171_/X vssd1 vssd1 vccd1 vccd1 _13979_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1787 _14661_/Q vssd1 vssd1 vccd1 vccd1 hold1787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1798 _11963_/X vssd1 vssd1 vccd1 vccd1 _14782_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07769_ _13674_/A1 hold1987/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15437_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11723__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ _10246_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12978__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09701__B _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12522__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10780_ _11580_/A _11578_/A _14968_/Q vssd1 vssd1 vccd1 vccd1 _10781_/B sky130_fd_sc_hd__and3_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09252_/X _09254_/X _09437_/Y _09438_/X vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08317__B _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _12446_/X _12447_/X _12449_/X _12448_/X _12644_/A1 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12451_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ _11401_/A _11401_/B vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__nor2_1
X_12381_ _13027_/A _12378_/X _12380_/X vssd1 vssd1 vccd1 vccd1 _13142_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_80 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_91 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07648__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14120_ _15191_/CLK _14120_/D vssd1 vssd1 vccd1 vccd1 _14120_/Q sky130_fd_sc_hd__dfxtp_1
X_11332_ _11333_/B _15223_/Q _15224_/Q _11526_/A vssd1 vssd1 vccd1 vccd1 _11334_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14051_ _15424_/CLK _14051_/D vssd1 vssd1 vccd1 vccd1 _14051_/Q sky130_fd_sc_hd__dfxtp_1
X_11263_ _11328_/A _11261_/X _11073_/Y _11076_/X vssd1 vssd1 vccd1 vccd1 _11264_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12589__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ _13102_/A _13002_/B _13002_/C vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__and3_1
X_10214_ _09970_/Y _09973_/Y _10392_/A _10213_/X vssd1 vssd1 vccd1 vccd1 _10392_/B
+ sky130_fd_sc_hd__a211oi_2
X_11194_ _11542_/A _11536_/A _11537_/B _11378_/C vssd1 vssd1 vccd1 vccd1 _11382_/A
+ sky130_fd_sc_hd__nand4_2
X_10145_ _10022_/A _10316_/B _10312_/A _10144_/D vssd1 vssd1 vccd1 vccd1 _10145_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09164__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _07261_/A _09915_/X _07319_/D vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__a21o_1
X_14953_ _14954_/CLK _14953_/D vssd1 vssd1 vccd1 vccd1 _14953_/Q sky130_fd_sc_hd__dfxtp_2
X_13904_ _15416_/CLK _13904_/D vssd1 vssd1 vccd1 vccd1 _13904_/Q sky130_fd_sc_hd__dfxtp_1
X_14884_ _14889_/CLK _14884_/D vssd1 vssd1 vccd1 vccd1 _14884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10772__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12418__A1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13835_ _14754_/CLK _13835_/D vssd1 vssd1 vccd1 vccd1 _13835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15045_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_203_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13414__A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ hold229/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10994_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07412__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _12917_/A1 _12716_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_169_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13697_ hold1843/X _13730_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 _13697_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15436_ _15436_/CLK _15436_/D vssd1 vssd1 vccd1 vccd1 _15436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ hold235/A _14311_/Q hold697/A _13971_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12648_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12456__A1_N _08107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15367_ _15367_/CLK hold340/X vssd1 vssd1 vccd1 vccd1 hold339/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _08532_/Y _12325_/B _12578_/X vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_170_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ _15376_/CLK _14318_/D vssd1 vssd1 vccd1 vccd1 _14318_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11588__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ _15301_/CLK _15298_/D vssd1 vssd1 vccd1 vccd1 _15298_/Q sky130_fd_sc_hd__dfxtp_1
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 hold328/A vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold339 hold339/A vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14249_ _15442_/CLK hold602/X vssd1 vssd1 vccd1 vccd1 hold601/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2349_A _15034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 _14489_/Q vssd1 vssd1 vccd1 vccd1 _12365_/S1 sky130_fd_sc_hd__buf_4
Xfanout819 _12460_/S vssd1 vssd1 vccd1 vccd1 _12491_/S sky130_fd_sc_hd__buf_6
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _08926_/A _09864_/A _08810_/C _08922_/A vssd1 vssd1 vccd1 vccd1 _08922_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__09770__A1 _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11808__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ hold447/A _15282_/Q _15090_/Q _14383_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09790_/X sky130_fd_sc_hd__mux4_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _11930_/X vssd1 vssd1 vccd1 vccd1 _14750_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _15088_/Q vssd1 vssd1 vccd1 vccd1 hold1017/X sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _08741_/A _09344_/B vssd1 vssd1 vccd1 vccd1 _08743_/C sky130_fd_sc_hd__and2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1028 _07481_/X vssd1 vssd1 vccd1 vccd1 _14109_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1039 _15069_/Q vssd1 vssd1 vccd1 vccd1 hold1039/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08672_ _09009_/A _09136_/A _09858_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _08673_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07306__B _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07623_ hold1819/X _13729_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07623_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10948__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15324_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07554_ _13386_/A hold131/X vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__and2_1
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09825__A2 _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07485_ hold1093/X _13724_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07836__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ hold223/A hold637/A _14606_/Q _13975_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09224_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09155_ _09154_/B _09154_/C _09154_/A vssd1 vssd1 vccd1 vccd1 _09157_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_A _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08106_ _08107_/A hold443/X vssd1 vssd1 vccd1 vccd1 _08106_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09086_ _09086_/A _09086_/B vssd1 vssd1 vccd1 vccd1 _13357_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ _08038_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__or2_1
XFILLER_0_13_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold840 hold840/A vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 hold851/A vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold862 hold862/A vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A1 _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold873 hold873/A vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 hold884/A vssd1 vssd1 vccd1 vccd1 hold884/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 hold895/A vssd1 vssd1 vccd1 vccd1 hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11718__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07998__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _09987_/B _09987_/C _09987_/A vssd1 vssd1 vccd1 vccd1 _09988_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2230 _07134_/X vssd1 vssd1 vccd1 vccd1 _13944_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2241 _14462_/Q vssd1 vssd1 vccd1 vccd1 hold2241/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2252 _11655_/X vssd1 vssd1 vccd1 vccd1 _14458_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08939_ _08940_/A _08940_/B _08940_/C vssd1 vssd1 vccd1 vccd1 _08939_/X sky130_fd_sc_hd__and3_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2263 _14728_/Q vssd1 vssd1 vccd1 vccd1 hold2263/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12122__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2274 _07092_/X vssd1 vssd1 vccd1 vccd1 _13905_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08316__A2 _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1540 _11880_/X vssd1 vssd1 vccd1 vccd1 _14702_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2285 _13926_/Q vssd1 vssd1 vccd1 vccd1 hold2285/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1551 _13813_/Q vssd1 vssd1 vccd1 vccd1 hold1551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2296 _13516_/X vssd1 vssd1 vccd1 vccd1 _15274_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11950_ _13705_/A1 hold1439/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11950_/X sky130_fd_sc_hd__mux2_1
Xhold1562 _07735_/X vssd1 vssd1 vccd1 vccd1 _14354_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1573 _14540_/Q vssd1 vssd1 vccd1 vccd1 hold1573/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1584 _11972_/X vssd1 vssd1 vccd1 vccd1 _14791_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _10900_/A _10900_/B _11089_/B _10900_/D vssd1 vssd1 vccd1 vccd1 _10901_/Y
+ sky130_fd_sc_hd__o22ai_2
Xhold1595 _14481_/Q vssd1 vssd1 vccd1 vccd1 hold1595/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ hold911/X _13735_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold912/A sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _07433_/A _13625_/C _13619_/X _13622_/C1 vssd1 vssd1 vccd1 vccd1 _15337_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ _10642_/X _10645_/X _10830_/Y _10831_/X vssd1 vssd1 vccd1 vccd1 _10832_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07232__A _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13551_ _08253_/B _08441_/B _13550_/X _13541_/A vssd1 vssd1 vccd1 vccd1 _13551_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ _11493_/A _10763_/B vssd1 vssd1 vccd1 vccd1 _10763_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _13027_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _13490_/A hold3/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__and2_1
XFILLER_0_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10694_ _10694_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15221_ _15225_/CLK _15221_/D vssd1 vssd1 vccd1 vccd1 _15221_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11689__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ hold1529/X hold2239/X hold1215/X hold1167/X _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12433_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11387__A1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__B2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15152_ _15304_/CLK _15152_/D vssd1 vssd1 vccd1 vccd1 _15152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ _12360_/X _12361_/X _12363_/X _12362_/X _12366_/A _06944_/A vssd1 vssd1 vccd1
+ vccd1 _12364_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08063__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10595__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14103_ _14105_/CLK hold244/X vssd1 vssd1 vccd1 vccd1 _14103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11315_ _11497_/A _11315_/B vssd1 vssd1 vccd1 vccd1 _11315_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15083_ _15372_/CLK _15083_/D vssd1 vssd1 vccd1 vccd1 _15083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12295_ _07438_/A _14087_/Q _14090_/Q _12294_/A vssd1 vssd1 vccd1 vccd1 _12295_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11139__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14034_ _15425_/CLK _14034_/D vssd1 vssd1 vccd1 vccd1 _14034_/Q sky130_fd_sc_hd__dfxtp_1
X_11246_ _11517_/A _15221_/Q _11247_/C _11348_/A vssd1 vssd1 vccd1 vccd1 _11248_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08004__B2 _13176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12887__A1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output253_A _14427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _11177_/A _11177_/B _11177_/C vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10128_ _10827_/C _10126_/X _10127_/X vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10059_ _10056_/Y _10057_/X _09896_/C _09896_/Y vssd1 vssd1 vccd1 vccd1 _10059_/X
+ sky130_fd_sc_hd__a211o_1
X_14936_ _15256_/CLK _14936_/D vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14867_ _14876_/CLK _14867_/D vssd1 vssd1 vccd1 vccd1 _14867_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12459__S _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__D _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13144__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818_ _15376_/CLK _13818_/D vssd1 vssd1 vccd1 vccd1 _13818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12498__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ _15188_/CLK _14798_/D vssd1 vssd1 vccd1 vccd1 _14798_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10487__B _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09363__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07818__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _13749_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13749_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12811__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ _11537_/B _09724_/D vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15419_ _15456_/CLK _15419_/D vssd1 vssd1 vccd1 vccd1 _15419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__buf_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10008__A _15200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15309_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _09911_/A _09911_/B vssd1 vssd1 vccd1 vccd1 _09911_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__buf_1
XFILLER_0_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12878__B2 _13194_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 _15209_/Q vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__clkbuf_4
Xfanout616 _08685_/C vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09842_ _09958_/B _09841_/C _09841_/A vssd1 vssd1 vccd1 vccd1 _09842_/Y sky130_fd_sc_hd__a21oi_2
Xfanout627 _15203_/Q vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__buf_6
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout638 _15200_/Q vssd1 vssd1 vccd1 vccd1 _08012_/B sky130_fd_sc_hd__clkbuf_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12973__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout649 _15198_/Q vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__buf_4
XANTENNA__12223__A _13374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07317__A _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _10744_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__or2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _13657_/A1 hold1357/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06985_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _08721_/Y _08722_/X _08617_/B _08617_/Y vssd1 vssd1 vccd1 vccd1 _08725_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__12725__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07751__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08989_/A _08652_/X _08654_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08656_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10678__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12369__S _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout549_A _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08793__D _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07606_ _13745_/A1 hold835/X _07609_/S vssd1 vssd1 vccd1 vccd1 hold836/A sky130_fd_sc_hd__mux2_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13055__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08586_ _08586_/A _08586_/B _08586_/C vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12489__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07537_ hold467/X _13708_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold468/A sky130_fd_sc_hd__mux2_1
XFILLER_0_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout716_A _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _13535_/B hold111/X vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__and2_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09207_ _12221_/B _09205_/Y _09340_/B _08526_/B hold2558/X vssd1 vssd1 vccd1 vccd1
+ _09207_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_106_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09106__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ _07852_/B _07475_/B vssd1 vssd1 vccd1 vccd1 _14029_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07198__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ _09138_/A _09712_/B _09138_/C _09138_/D vssd1 vssd1 vccd1 vccd1 _09138_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_115_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ _09199_/B _09069_/B vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_60_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ _10959_/X _10960_/X _11099_/Y vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__12869__A1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _14980_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12080_/X
+ sky130_fd_sc_hd__or4_1
Xhold670 hold670/A vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10860__B _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 hold681/A vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 hold692/A vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _10847_/X _10850_/X _11029_/X _11030_/Y vssd1 vssd1 vccd1 vccd1 _11033_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09426__B _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2060 _07094_/X vssd1 vssd1 vccd1 vccd1 _13907_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2071 _13809_/Q vssd1 vssd1 vccd1 vccd1 hold2071/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13663__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2082 _07095_/X vssd1 vssd1 vccd1 vccd1 _13908_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13294__A1 input137/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _13107_/A _12982_/B vssd1 vssd1 vccd1 vccd1 _14967_/D sky130_fd_sc_hd__nor2_1
Xhold2093 _14208_/Q vssd1 vssd1 vccd1 vccd1 hold2093/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07661__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1370 _07734_/X vssd1 vssd1 vccd1 vccd1 _14353_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1381 _13883_/Q vssd1 vssd1 vccd1 vccd1 hold1381/X sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ _15265_/CLK _14721_/D vssd1 vssd1 vccd1 vccd1 _14721_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _13655_/A1 hold1881/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11933_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1392 _07620_/X vssd1 vssd1 vccd1 vccd1 _14243_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _15387_/CLK hold788/X vssd1 vssd1 vccd1 vccd1 hold787/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11864_ hold343/X _13718_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold344/A sky130_fd_sc_hd__mux2_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13603_ _07424_/A _13625_/C _13602_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15328_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10814_/B _10814_/C _10814_/A vssd1 vssd1 vccd1 vccd1 _10817_/C sky130_fd_sc_hd__a21o_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _15416_/CLK hold242/X vssd1 vssd1 vccd1 vccd1 hold241/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ hold557/X _13748_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold558/A sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11911__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _15068_/Q hold769/X _13534_/S vssd1 vssd1 vccd1 vccd1 hold770/A sky130_fd_sc_hd__mux2_1
XFILLER_0_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10746_ _10746_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _11108_/C sky130_fd_sc_hd__or2_1
XFILLER_0_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _11291_/B _13468_/A _13464_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 _13465_/X
+ sky130_fd_sc_hd__o211a_1
X_10677_ _10677_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10717_/A sky130_fd_sc_hd__or2_1
XFILLER_0_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15204_ _15324_/CLK _15204_/D vssd1 vssd1 vccd1 vccd1 _15204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09648__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12416_ hold603/A _14238_/Q _12459_/S vssd1 vssd1 vccd1 vccd1 _12416_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13396_ _13396_/A _13396_/B vssd1 vssd1 vccd1 vccd1 _15187_/D sky130_fd_sc_hd__and2_1
XFILLER_0_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10032__A1 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__B2 _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__D _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput208 _14190_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[20] sky130_fd_sc_hd__buf_12
XFILLER_0_65_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15135_ _15320_/CLK _15135_/D vssd1 vssd1 vccd1 vccd1 _15135_/Q sky130_fd_sc_hd__dfxtp_1
X_12347_ _14782_/Q _14494_/Q _12466_/S vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__mux2_1
Xoutput219 _14200_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[30] sky130_fd_sc_hd__buf_12
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ _15068_/CLK _15066_/D vssd1 vssd1 vccd1 vccd1 _15066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12278_ _13389_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _14927_/D sky130_fd_sc_hd__nor2_2
XANTENNA__09725__A1 _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ _15385_/CLK hold776/X vssd1 vssd1 vccd1 vccd1 hold775/A sky130_fd_sc_hd__dfxtp_1
X_11229_ _11229_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11231_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07831__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13285__A1 input134/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09352__A _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__B1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ _15244_/CLK _14919_/D vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__A2 _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _08440_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08440_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13037__A1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08873_/A _08370_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _08371_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10010__B _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11821__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ _10600_/B _09075_/B _10951_/B vssd1 vssd1 vccd1 vccd1 _07330_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08464__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2750_A _15173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07253_ _15224_/Q _14968_/Q vssd1 vssd1 vccd1 vccd1 _07253_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07184_ hold1647/X _13652_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07184_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13748__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07746__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__B _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _07477_/Y vssd1 vssd1 vccd1 vccd1 _07509_/S sky130_fd_sc_hd__clkbuf_16
Xfanout413 _06978_/X vssd1 vssd1 vccd1 vccd1 _06994_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__09246__B _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12946__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 _11961_/Y vssd1 vssd1 vccd1 vccd1 _11993_/S sky130_fd_sc_hd__buf_12
Xfanout435 _07710_/X vssd1 vssd1 vccd1 vccd1 _07726_/S sky130_fd_sc_hd__clkbuf_16
Xfanout446 hold2520/X vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__clkbuf_4
X_09825_ _09979_/B _11588_/A _11623_/A _10183_/A vssd1 vssd1 vccd1 vccd1 _09828_/C
+ sky130_fd_sc_hd__a22o_1
Xfanout457 _12195_/A2 vssd1 vssd1 vccd1 vccd1 _12173_/A2 sky130_fd_sc_hd__buf_4
Xfanout468 _07884_/X vssd1 vssd1 vccd1 vccd1 _12258_/S sky130_fd_sc_hd__buf_8
Xfanout479 _06959_/X vssd1 vssd1 vccd1 vccd1 _10949_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout666_A _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09756_ _09608_/X _09610_/Y _09754_/X _09755_/Y vssd1 vssd1 vccd1 vccd1 _09910_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13276__A1 input131/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ _14082_/Q _14081_/Q _06968_/C vssd1 vssd1 vccd1 vccd1 _06972_/C sky130_fd_sc_hd__or3_1
XANTENNA__07481__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _08707_/A _08805_/A _08707_/C vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09262__A _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09687_ _09683_/X _09685_/Y _09547_/B _09549_/B vssd1 vssd1 vccd1 vccd1 _09687_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout833_A _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08638_ _08964_/B _07912_/X _08637_/Y vssd1 vssd1 vccd1 vccd1 _08640_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13028__B2 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08569_ _08569_/A _08569_/B _08569_/C vssd1 vssd1 vccd1 vccd1 _08569_/X sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_4_0__f_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11731__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _10600_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ _11580_/A _14972_/Q vssd1 vssd1 vccd1 vccd1 _11581_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _10696_/B _10530_/C _10530_/A vssd1 vssd1 vccd1 vccd1 _10532_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12128__A _12128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ input87/X fanout1/X _13249_/X vssd1 vssd1 vccd1 vccd1 _13251_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08207__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ _10463_/A _10463_/B _10463_/C vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11389__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13658__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _12247_/A _12196_/X _12200_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _12208_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09955__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13751__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ _13481_/A _13181_/B vssd1 vssd1 vccd1 vccd1 _15046_/D sky130_fd_sc_hd__and2_1
X_10393_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07656__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09437__A _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _14877_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09707__A1 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _12063_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _14844_/D sky130_fd_sc_hd__and2_1
XANTENNA__09707__B2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08066__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__B1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__B2 _13203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11014_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_198_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07813__S0 _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13267__A1 input159/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ hold2213/X hold1007/X _13066_/S vssd1 vssd1 vccd1 vccd1 _12965_/X sky130_fd_sc_hd__mux2_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08143__B1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _13671_/A1 hold1737/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__mux2_1
X_14704_ _15446_/CLK _14704_/D vssd1 vssd1 vccd1 vccd1 _14704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__A1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _15381_/Q _15284_/Q _15092_/Q _14385_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12896_/X sky130_fd_sc_hd__mux4_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14731_/CLK hold888/X vssd1 vssd1 vccd1 vccd1 hold887/A sky130_fd_sc_hd__dfxtp_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ hold1059/X _13734_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__mux2_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12778__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _15270_/CLK hold226/X vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__dfxtp_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ hold1589/X _13665_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11778_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12873__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13141__B _13141_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ _13665_/A1 hold1283/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10729_ _10728_/B _10728_/C _10728_/A vssd1 vssd1 vccd1 vccd1 _10730_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14497_ _15265_/CLK hold484/X vssd1 vssd1 vccd1 vccd1 hold483/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13448_ _13450_/A _13448_/B vssd1 vssd1 vccd1 vccd1 _13448_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12625__S0 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_173_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10781__A _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ _13386_/A _13379_/B vssd1 vssd1 vccd1 vccd1 _15170_/D sky130_fd_sc_hd__and2_1
X_15118_ _15127_/CLK _15118_/D vssd1 vssd1 vccd1 vccd1 _15118_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_53_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__B _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold2331_A _15342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _08201_/A _07940_/B vssd1 vssd1 vccd1 vccd1 _07940_/Y sky130_fd_sc_hd__nor2_1
X_15049_ _15440_/CLK _15049_/D vssd1 vssd1 vccd1 vccd1 _15049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_11__f_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2807 _12744_/X vssd1 vssd1 vccd1 vccd1 _12745_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13050__S0 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_188_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2818 _14221_/Q vssd1 vssd1 vccd1 vccd1 hold2818/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2829 _15323_/Q vssd1 vssd1 vccd1 vccd1 hold2829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07871_ _07862_/B _14087_/Q _07744_/A _15343_/Q vssd1 vssd1 vccd1 vccd1 _07871_/X
+ sky130_fd_sc_hd__a22o_1
X_09610_ _09394_/X _09397_/X _09608_/X _09609_/Y vssd1 vssd1 vccd1 vccd1 _09610_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_177_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11816__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13258__A1 input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09541_ _09979_/B _15209_/Q _09860_/B _10183_/A vssd1 vssd1 vccd1 vccd1 _09543_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_111_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15234__D _15234_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09472_ _09471_/B _09471_/C _09471_/A vssd1 vssd1 vccd1 vccd1 _09472_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07314__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08423_ _08519_/A _08421_/Y _08317_/C _08318_/C vssd1 vssd1 vccd1 vccd1 _08427_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_126_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ _08544_/C _08353_/Y _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_163_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12864__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07305_ _08569_/B _07305_/B vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ _12252_/B _08285_/B vssd1 vssd1 vccd1 vccd1 _08285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_172_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout414_A _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ _08075_/B _11566_/A vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09937__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _13668_/A1 hold1627/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07167_/X sky130_fd_sc_hd__mux2_1
X_07098_ _13734_/A1 hold1793/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07098_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout783_A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11726__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _10338_/B _09809_/C _11536_/B _10166_/A vssd1 vssd1 vccd1 vccd1 _09808_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__13249__A1 input151/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _09739_/A _09739_/B _09739_/C vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__and3_1
XFILLER_0_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12750_ _12746_/X _12747_/X _12749_/X _12748_/X _12844_/A1 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12751_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_167_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11701_ hold483/X _13655_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold484/A sky130_fd_sc_hd__mux2_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11680__A0 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12681_ _13106_/A1 _13154_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__o21a_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14775_/CLK _14420_/D vssd1 vssd1 vccd1 vccd1 _14420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11632_ _11632_/A _11632_/B vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__xnor2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10235__A1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _15090_/CLK hold384/X vssd1 vssd1 vccd1 vccd1 hold383/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ _11563_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _13317_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _15120_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_123_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11983__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ _10513_/A _10513_/B _10513_/C vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14282_ _14472_/CLK _14282_/D vssd1 vssd1 vccd1 vccd1 _14282_/Q sky130_fd_sc_hd__dfxtp_1
X_11494_ _14297_/Q _14233_/Q _14169_/Q _14487_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11495_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13233_ hold411/X _13679_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold412/A sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _13390_/A _13164_/B vssd1 vssd1 vccd1 vccd1 _15029_/D sky130_fd_sc_hd__nor2_1
X_10376_ _10372_/Y _10374_/X _10156_/X _10160_/B vssd1 vssd1 vccd1 vccd1 _10376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output166_A _15178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ hold2459/X _12129_/A2 _12114_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12115_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13095_ _13095_/A _13095_/B _13076_/A vssd1 vssd1 vccd1 vccd1 _13102_/B sky130_fd_sc_hd__or3b_1
X_12046_ _12112_/A hold2698/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12047_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09787__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__B1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output333_A _14831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13997_ _15365_/CLK hold718/X vssd1 vssd1 vccd1 vccd1 hold717/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ hold163/A hold627/A hold485/A _13983_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12948_/X sky130_fd_sc_hd__mux4_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11671__A0 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_170 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ _13396_/B _13104_/A2 _12878_/X vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10776__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__S0 _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13152__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_181 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_192 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _15421_/CLK _14618_/D vssd1 vssd1 vccd1 vccd1 _14618_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12846__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14549_ _15451_/CLK _14549_/D vssd1 vssd1 vccd1 vccd1 _14549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09092__A1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08070_ _12252_/B _08070_/B vssd1 vssd1 vccd1 vccd1 _08070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_113_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07021_ hold905/X _13659_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 hold906/A sky130_fd_sc_hd__mux2_1
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10529__A2 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09077__A _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08972_ _09494_/A1 _08862_/Y _08971_/X vssd1 vssd1 vccd1 vccd1 _08972_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13023__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2604 _15331_/Q vssd1 vssd1 vccd1 vccd1 _07353_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2615 _14439_/Q vssd1 vssd1 vccd1 vccd1 _09087_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2626 _12155_/X vssd1 vssd1 vccd1 vccd1 _14888_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _14426_/Q _13586_/B vssd1 vssd1 vccd1 vccd1 _07923_/Y sky130_fd_sc_hd__nor2_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2637 _14889_/Q vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2648 _15105_/Q vssd1 vssd1 vccd1 vccd1 hold2648/X sky130_fd_sc_hd__buf_1
XANTENNA__12151__A1 hold2607/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1903 _14743_/Q vssd1 vssd1 vccd1 vccd1 hold1903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2659 _14820_/Q vssd1 vssd1 vccd1 vccd1 hold2659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1914 _07075_/X vssd1 vssd1 vccd1 vccd1 _13891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1925 _14248_/Q vssd1 vssd1 vccd1 vccd1 hold1925/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09524__B _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ _07855_/A _07857_/C _07855_/C vssd1 vssd1 vccd1 vccd1 _07854_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1936 _06987_/X vssd1 vssd1 vccd1 vccd1 _13806_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1947 _15449_/Q vssd1 vssd1 vccd1 vccd1 hold1947/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12231__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10701__A2 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1958 _07144_/X vssd1 vssd1 vccd1 vccd1 _13954_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1969 _13830_/Q vssd1 vssd1 vccd1 vccd1 hold1969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07785_ hold1735/X _13690_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 _07785_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09524_ _09661_/A _09809_/C vssd1 vssd1 vccd1 vccd1 _09527_/A sky130_fd_sc_hd__and2_1
XFILLER_0_211_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08202__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09270_/Y _09273_/X _09453_/Y _09454_/X vssd1 vssd1 vccd1 vccd1 _09557_/A
+ sky130_fd_sc_hd__a211oi_4
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08753__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07979__B _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout629_A _15202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _08406_/A _08406_/B vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_136_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09386_ _10166_/A _10338_/B _09676_/D _09979_/C vssd1 vssd1 vccd1 vccd1 _09387_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08337_ _10397_/A _08380_/B _08337_/C vssd1 vssd1 vccd1 vccd1 _08337_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_35_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07995__A _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ _08877_/A _08267_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08268_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07219_ _14066_/Q _14065_/Q vssd1 vssd1 vccd1 vccd1 _07856_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08199_ _08201_/A _08199_/B vssd1 vssd1 vccd1 vccd1 _08199_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08603__B _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ _10401_/C _10230_/B vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11193__A2 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _10160_/B _10160_/C _10160_/A vssd1 vssd1 vccd1 vccd1 _10164_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__12840__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10092_ _10244_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_195_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13237__A _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13920_ _15453_/CLK _13920_/D vssd1 vssd1 vccd1 vccd1 _13920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13851_ _15089_/CLK hold398/X vssd1 vssd1 vccd1 vccd1 hold397/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09153__C _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ _13102_/A _12802_/B _12802_/C vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13782_ hold241/X vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10994_ _10994_/A _10994_/B _10994_/C vssd1 vssd1 vccd1 vccd1 _10996_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_96_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _15407_/Q hold693/A _14702_/Q _14766_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12733_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07889__B _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15452_/CLK hold438/X vssd1 vssd1 vccd1 vccd1 hold437/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ hold799/X hold2798/X hold701/X hold1555/X _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12664_/X sky130_fd_sc_hd__mux4_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14403_ _15045_/CLK hold926/X vssd1 vssd1 vccd1 vccd1 hold925/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11615_ _11567_/A _15227_/Q _11346_/A _11344_/A vssd1 vssd1 vccd1 vccd1 _11617_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_182_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__B _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15383_ _15383_/CLK _15383_/D vssd1 vssd1 vccd1 vccd1 _15383_/Q sky130_fd_sc_hd__dfxtp_1
X_12595_ _12595_/A _12595_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _15042_/CLK hold604/X vssd1 vssd1 vccd1 vccd1 hold603/A sky130_fd_sc_hd__dfxtp_1
X_11546_ _11546_/A _11546_/B vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ _15456_/CLK _14265_/D vssd1 vssd1 vccd1 vccd1 _14265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11477_ _11645_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11479_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ hold981/X _13662_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 hold982/A sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10428_ _11504_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10428_/Y sky130_fd_sc_hd__nor2_1
X_14196_ _15188_/CLK _14196_/D vssd1 vssd1 vccd1 vccd1 _14196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12381__A1 _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13381_/A _13147_/B vssd1 vssd1 vccd1 vccd1 _15012_/D sky130_fd_sc_hd__nor2_1
X_10359_ _11517_/A _10166_/C _10524_/A _10358_/D vssd1 vssd1 vccd1 vccd1 _10360_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12669__C1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13078_ _13714_/A1 _13103_/A2 _13078_/B1 _13202_/B vssd1 vssd1 vccd1 vccd1 _13078_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12133__A1 _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12029_ _12063_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _14827_/D sky130_fd_sc_hd__and2_1
XANTENNA__13147__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07570_ _13397_/A hold167/X vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__and2_1
XANTENNA__13094__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__C _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12197__S _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09240_ _09941_/A _09239_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09240_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09171_ _10185_/A _09858_/C _09171_/C _09297_/A vssd1 vssd1 vccd1 vccd1 _09297_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08122_ _08201_/A _08119_/X _08121_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _08123_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08273__C1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _08201_/A _08052_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08053_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_82_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07004_ _11921_/A0 hold761/X _07010_/S vssd1 vssd1 vccd1 vccd1 hold762/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07379__A1 _15341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08142__C _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12660__S _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2401 _13563_/X vssd1 vssd1 vccd1 vccd1 _15307_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07754__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput108 in1[1] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__clkbuf_1
X_08955_ _08955_/A _08955_/B vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__xnor2_2
Xhold2412 _14068_/Q vssd1 vssd1 vccd1 vccd1 _07410_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput119 in1[2] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_1
Xhold2423 _12091_/X vssd1 vssd1 vccd1 vccd1 _14857_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2434 _12079_/X vssd1 vssd1 vccd1 vccd1 _14851_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout579_A _15220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1700 _07102_/X vssd1 vssd1 vccd1 vccd1 _13915_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2445 _13461_/X vssd1 vssd1 vccd1 vccd1 _15224_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _13241_/A _07910_/B _07904_/B vssd1 vssd1 vccd1 vccd1 _07908_/C sky130_fd_sc_hd__or3b_1
Xhold1711 _13932_/Q vssd1 vssd1 vccd1 vccd1 hold1711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2456 _12109_/X vssd1 vssd1 vccd1 vccd1 _14866_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08886_ _09571_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__nand2_1
Xhold2467 _14868_/Q vssd1 vssd1 vccd1 vccd1 hold2467/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08879__A1 _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1722 _07141_/X vssd1 vssd1 vccd1 vccd1 _13951_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1733 _13930_/Q vssd1 vssd1 vccd1 vccd1 hold1733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2478 _09925_/X vssd1 vssd1 vccd1 vccd1 hold2478/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2489 _14873_/Q vssd1 vssd1 vccd1 vccd1 hold2489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07000__A0 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1744 _07104_/X vssd1 vssd1 vccd1 vccd1 _13917_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1755 _14698_/Q vssd1 vssd1 vccd1 vccd1 hold1755/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09540__A2 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07837_ _14028_/Q _14029_/Q _06950_/X _06959_/X vssd1 vssd1 vccd1 vccd1 _12308_/B
+ sky130_fd_sc_hd__o31ai_2
Xhold1766 _13713_/X vssd1 vssd1 vccd1 vccd1 _15419_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1777 _14477_/Q vssd1 vssd1 vccd1 vccd1 hold1777/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_A _14953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1788 _11838_/X vssd1 vssd1 vccd1 vccd1 _14661_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1799 _14764_/Q vssd1 vssd1 vccd1 vccd1 hold1799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07768_ _13673_/A1 hold2041/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07768_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10438__A1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _09514_/A _09504_/X _09506_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09508_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09701__C _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ hold1649/X _13738_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 _07699_/X sky130_fd_sc_hd__mux2_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09714_/A _09712_/B _09437_/C _09437_/D vssd1 vssd1 vccd1 vccd1 _09438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09369_ hold673/A _14220_/Q hold305/A hold587/A _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09370_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_118_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12835__S _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _11399_/B _11399_/C _11399_/A vssd1 vssd1 vccd1 vccd1 _11401_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12060__A0 hold2610/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12380_ _13174_/B _12953_/B1 _12354_/X _13653_/A1 _12379_/X vssd1 vssd1 vccd1 vccd1
+ _12380_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_117_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_70 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_81 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10610__A1 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_92 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10610__B2 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12136__A _14879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11040__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14050_ _14083_/CLK hold196/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_11262_ _11073_/Y _11076_/X _11328_/A _11261_/X vssd1 vssd1 vccd1 vccd1 _11328_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _13101_/A _13001_/B vssd1 vssd1 vccd1 vccd1 _13002_/C sky130_fd_sc_hd__or2_1
X_10213_ _10386_/B _10211_/X _10058_/Y _10060_/Y vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13666__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _11536_/A _11537_/B _11378_/C _11542_/A vssd1 vssd1 vccd1 vccd1 _11196_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07664__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10144_ _11563_/A _10316_/B _10312_/A _10144_/D vssd1 vssd1 vccd1 vccd1 _10312_/B
+ sky130_fd_sc_hd__nand4_2
Xclkbuf_2_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09164__B _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ _10397_/A _10075_/B _10220_/B vssd1 vssd1 vccd1 vccd1 _10075_/X sky130_fd_sc_hd__or3_2
X_14952_ _15222_/CLK _14952_/D vssd1 vssd1 vccd1 vccd1 _14952_/Q sky130_fd_sc_hd__dfxtp_1
X_13903_ _15436_/CLK _13903_/D vssd1 vssd1 vccd1 vccd1 _13903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14883_ _14889_/CLK _14883_/D vssd1 vssd1 vccd1 vccd1 _14883_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07542__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11914__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13834_ _14595_/CLK hold810/X vssd1 vssd1 vccd1 vccd1 hold809/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13765_ hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10977_ _10976_/A _10976_/B _10791_/Y vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_202_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07412__B _07412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12716_ hold539/A hold545/A _12791_/S vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13696_ hold803/X _13729_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 hold804/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ hold785/A hold725/A _14634_/Q _14730_/Q _12641_/S _12689_/S1 vssd1 vssd1
+ vccd1 vccd1 _12647_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ _15435_/CLK _15435_/D vssd1 vssd1 vccd1 vccd1 _15435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15366_ _15400_/CLK _15366_/D vssd1 vssd1 vccd1 vccd1 _15366_/Q sky130_fd_sc_hd__dfxtp_1
X_12578_ _13661_/A1 _12329_/B _12953_/B1 _13182_/B vssd1 vssd1 vccd1 vccd1 _12578_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11555_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14317_ _15372_/CLK hold538/X vssd1 vssd1 vccd1 vccd1 hold537/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15297_ _15320_/CLK _15297_/D vssd1 vssd1 vccd1 vccd1 _15297_/Q sky130_fd_sc_hd__dfxtp_1
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 hold329/A vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ _15191_/CLK _14248_/D vssd1 vssd1 vccd1 vccd1 _14248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _15177_/CLK hold132/X vssd1 vssd1 vccd1 vccd1 _14179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08653__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 _12899_/S1 vssd1 vssd1 vccd1 vccd1 _12749_/S1 sky130_fd_sc_hd__clkbuf_8
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__C1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ _09344_/B _10744_/A vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__and2b_4
Xhold1007 _14132_/Q vssd1 vssd1 vccd1 vccd1 hold1007/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _13224_/X vssd1 vssd1 vccd1 vccd1 _15088_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold2509_A _14988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1029 _13836_/Q vssd1 vssd1 vccd1 vccd1 hold1029/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08671_ _08776_/A _09858_/A _09858_/B _09009_/A vssd1 vssd1 vccd1 vccd1 _08673_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_205_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11824__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ hold973/X _13728_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 hold974/A sky130_fd_sc_hd__mux2_1
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2780_A _11287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07553_ _13393_/A hold151/X vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__and2_1
XFILLER_0_193_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11125__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ hold1531/X _13690_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09223_ _13570_/B _09221_/Y _09222_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _09223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12042__A0 hold2605/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _09154_/A _09154_/B _09154_/C vssd1 vssd1 vccd1 vccd1 _09157_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_161_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08434__A _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12593__A1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08105_ _08040_/A _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _08967_/B _08969_/B _08965_/X vssd1 vssd1 vccd1 vccd1 _09086_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_142_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08036_ _06903_/A _07433_/A _08036_/S vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__mux2_2
Xinput90 in0[3] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold830 hold830/A vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold841 hold841/A vssd1 vssd1 vccd1 vccd1 hold841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 hold852/A vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08549__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08013__A2 _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09210__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__S _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 hold863/A vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 hold874/A vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 hold885/A vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07484__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 hold896/A vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _09987_/A _09987_/B _09987_/C vssd1 vssd1 vccd1 vccd1 _09987_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_110_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2220 _11899_/X vssd1 vssd1 vccd1 vccd1 _14720_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout863_A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2231 _13940_/Q vssd1 vssd1 vccd1 vccd1 hold2231/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ _08935_/X _08936_/Y _08817_/Y _08819_/X vssd1 vssd1 vccd1 vccd1 _08940_/C
+ sky130_fd_sc_hd__a211o_1
Xhold2242 _11659_/X vssd1 vssd1 vccd1 vccd1 _14462_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2253 _14749_/Q vssd1 vssd1 vccd1 vccd1 hold2253/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2264 _11907_/X vssd1 vssd1 vccd1 vccd1 _14728_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1530 _13689_/X vssd1 vssd1 vccd1 vccd1 _15395_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2275 _14911_/Q vssd1 vssd1 vccd1 vccd1 _13472_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1541 _15083_/Q vssd1 vssd1 vccd1 vccd1 hold1541/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2286 _07116_/X vssd1 vssd1 vccd1 vccd1 _13926_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1552 _06994_/X vssd1 vssd1 vccd1 vccd1 _13813_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08869_/X sky130_fd_sc_hd__or2_1
Xhold2297 _13888_/Q vssd1 vssd1 vccd1 vccd1 hold2297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1563 _13898_/Q vssd1 vssd1 vccd1 vccd1 hold1563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1574 _11746_/X vssd1 vssd1 vccd1 vccd1 _14540_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _10900_/A _10900_/B _11089_/B _10900_/D vssd1 vssd1 vccd1 vccd1 _11085_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__11734__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1585 _14726_/Q vssd1 vssd1 vccd1 vccd1 hold1585/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ hold1539/X _13734_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__mux2_1
Xhold1596 _11678_/X vssd1 vssd1 vccd1 vccd1 _14481_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10831_ _11564_/A _10830_/B _10830_/C _10830_/D vssd1 vssd1 vccd1 vccd1 _10831_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07232__B _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ _14431_/Q _13554_/B vssd1 vssd1 vccd1 vccd1 _13550_/X sky130_fd_sc_hd__or2_1
X_10762_ hold563/A hold849/A hold481/A _14744_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10763_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _12676_/A _12501_/B vssd1 vssd1 vccd1 vccd1 _12502_/C sky130_fd_sc_hd__or2_1
XFILLER_0_164_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10831__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ _13481_/A _13481_/B vssd1 vssd1 vccd1 vccd1 _13481_/X sky130_fd_sc_hd__and2_1
X_10693_ _10873_/A _15223_/Q _10694_/A vssd1 vssd1 vccd1 vccd1 _10693_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12565__S _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15220_ _15222_/CLK _15220_/D vssd1 vssd1 vccd1 vccd1 _15220_/Q sky130_fd_sc_hd__dfxtp_2
X_12432_ _12482_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _14945_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08344__A _08345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11387__A2 _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15151_ _15304_/CLK _15151_/D vssd1 vssd1 vccd1 vccd1 _15151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _15392_/Q _14527_/Q _14687_/Q _14751_/Q _12365_/S0 _12343_/A vssd1 vssd1
+ vccd1 vccd1 _12363_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14102_ _14105_/CLK hold222/X vssd1 vssd1 vccd1 vccd1 _14102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11314_ hold487/A _13956_/Q hold399/A _13924_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _11315_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15082_ _15371_/CLK hold928/X vssd1 vssd1 vccd1 vccd1 hold927/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ _12294_/A _13241_/C _13240_/C vssd1 vssd1 vccd1 vccd1 _12294_/X sky130_fd_sc_hd__and3_1
XFILLER_0_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _15199_/CLK _14033_/D vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11909__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ _11541_/A _11351_/B _11586_/B _11620_/B vssd1 vssd1 vccd1 vccd1 _11348_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08004__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11544__C1 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _11173_/Y _11174_/X _10987_/D _10987_/Y vssd1 vssd1 vccd1 vccd1 _11177_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__B1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10127_ _10126_/B _11606_/A _10827_/C _10126_/A vssd1 vssd1 vccd1 vccd1 _10127_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10058_ _09896_/C _09896_/Y _10056_/Y _10057_/X vssd1 vssd1 vccd1 vccd1 _10058_/Y
+ sky130_fd_sc_hd__o211ai_4
X_14935_ _15256_/CLK _14935_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14866_ _14866_/CLK _14866_/D vssd1 vssd1 vccd1 vccd1 _14866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13144__B _13144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817_ _15439_/CLK _13817_/D vssd1 vssd1 vccd1 vccd1 _13817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14797_ _15374_/CLK _14797_/D vssd1 vssd1 vccd1 vccd1 _14797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09363__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ hold361/X _13748_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold362/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10784__A _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ hold1601/X _13679_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 _13679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12024__A0 _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15418_ _15418_/CLK hold808/X vssd1 vssd1 vccd1 vccd1 hold807/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15349_ _15425_/CLK _15349_/D vssd1 vssd1 vccd1 vccd1 _15349_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08874__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10008__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11819__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__nor2_1
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12422__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12878__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 _15209_/Q vssd1 vssd1 vccd1 vccd1 _09709_/B sky130_fd_sc_hd__buf_6
XFILLER_0_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09841_ _09841_/A _09958_/B _09841_/C vssd1 vssd1 vccd1 vccd1 _09841_/X sky130_fd_sc_hd__and3_2
Xfanout617 _15205_/Q vssd1 vssd1 vccd1 vccd1 _08685_/C sky130_fd_sc_hd__buf_4
Xfanout628 _15202_/Q vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__clkbuf_8
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout639 _11596_/A vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__buf_4
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07317__B _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _10744_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__nand2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _13656_/A1 hold1689/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06984_/X sky130_fd_sc_hd__mux2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08617_/B _08617_/Y _08721_/Y _08722_/X vssd1 vssd1 vccd1 vccd1 _08725_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13335__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08654_ _08981_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _08654_/X sky130_fd_sc_hd__or2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10678__B _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _13711_/A1 hold1597/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07605_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08585_ _08908_/A _09026_/B _09437_/A _08685_/C vssd1 vssd1 vccd1 vccd1 _08586_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout444_A _07389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12489__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07536_ hold645/X _13740_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold646/A sky130_fd_sc_hd__mux2_1
XFILLER_0_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07467_ _13501_/A hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__and2_1
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12385__S _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09206_ _09205_/B _09205_/C _09205_/A vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07479__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09106__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07398_ _07852_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14028_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09137_ _09138_/A _09712_/B _09138_/C _09138_/D vssd1 vssd1 vccd1 vccd1 _09137_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__A1 _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _09065_/A _09066_/X _08916_/X _08919_/X vssd1 vssd1 vccd1 vccd1 _09069_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08019_ _07961_/A _07961_/B _07959_/A vssd1 vssd1 vccd1 vccd1 _08020_/C sky130_fd_sc_hd__o21ai_1
Xhold660 hold660/A vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold671 hold671/A vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10860__C _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _11027_/Y _11028_/X _10814_/B _10817_/B vssd1 vssd1 vccd1 vccd1 _11030_/Y
+ sky130_fd_sc_hd__o211ai_4
Xhold682 hold682/A vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 hold693/A vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09426__C _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2050 _07048_/X vssd1 vssd1 vccd1 vccd1 _13864_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2061 _14739_/Q vssd1 vssd1 vccd1 vccd1 hold2061/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2072 _06990_/X vssd1 vssd1 vccd1 vccd1 _13809_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _13106_/A1 _12980_/Y _08637_/Y vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__o21a_1
Xhold2083 _13945_/Q vssd1 vssd1 vccd1 vccd1 hold2083/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2094 _07584_/X vssd1 vssd1 vccd1 vccd1 _14208_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1360 _07748_/X vssd1 vssd1 vccd1 vccd1 _14364_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13245__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _15264_/CLK _14720_/D vssd1 vssd1 vccd1 vccd1 _14720_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1371 _14376_/Q vssd1 vssd1 vccd1 vccd1 hold1371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1382 _07067_/X vssd1 vssd1 vccd1 vccd1 _13883_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ _13654_/A1 hold1309/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11932_/X sky130_fd_sc_hd__mux2_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1393 _14486_/Q vssd1 vssd1 vccd1 vccd1 hold1393/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14651_ _14651_/CLK hold342/X vssd1 vssd1 vccd1 vccd1 hold341/A sky130_fd_sc_hd__dfxtp_1
X_11863_ hold1379/X _12329_/A _11877_/S vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__mux2_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11057__A1 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10814_ _10814_/A _10814_/B _10814_/C vssd1 vssd1 vccd1 vccd1 _10817_/B sky130_fd_sc_hd__nand3_4
X_13602_ input55/X _13634_/B vssd1 vssd1 vccd1 vccd1 _13602_/X sky130_fd_sc_hd__or2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14582_ _15242_/CLK hold164/X vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__dfxtp_1
X_11794_ hold353/X _13681_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13533_ _13681_/A1 hold677/X _13534_/S vssd1 vssd1 vccd1 vccd1 hold678/A sky130_fd_sc_hd__mux2_1
X_10745_ _10745_/A _10745_/B vssd1 vssd1 vccd1 vccd1 _11108_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12006__A0 hold2586/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13464_ _13466_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13464_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08074__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _10673_/Y _10674_/X _10502_/B _10502_/Y vssd1 vssd1 vccd1 vccd1 _10676_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15203_ _15324_/CLK _15203_/D vssd1 vssd1 vccd1 vccd1 _15203_/Q sky130_fd_sc_hd__dfxtp_1
X_12415_ hold779/A _14110_/Q _12460_/S vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13395_ _13396_/A _13395_/B vssd1 vssd1 vccd1 vccd1 _15186_/D sky130_fd_sc_hd__and2_1
XFILLER_0_211_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10032__A2 _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15134_ _15460_/CLK _15134_/D vssd1 vssd1 vccd1 vccd1 _15134_/Q sky130_fd_sc_hd__dfxtp_1
X_12346_ hold883/A _15262_/Q _15070_/Q _14363_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12346_/X sky130_fd_sc_hd__mux4_1
Xoutput209 _14191_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[21] sky130_fd_sc_hd__buf_12
XFILLER_0_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ _15196_/CLK _15065_/D vssd1 vssd1 vccd1 vccd1 _15065_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09617__B _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ _13487_/A _12277_/B vssd1 vssd1 vccd1 vccd1 _14926_/D sky130_fd_sc_hd__and2_1
XANTENNA__12324__A _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ _14791_/CLK _14016_/D vssd1 vssd1 vccd1 vccd1 _14016_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09725__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _11228_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11231_/A sky130_fd_sc_hd__or2_1
XANTENNA__10415__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11159_ _11158_/B _11158_/C _11158_/A vssd1 vssd1 vccd1 vccd1 _11160_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10740__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13155__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14918_ _15196_/CLK _14918_/D vssd1 vssd1 vccd1 vccd1 _14918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14849_ _15254_/CLK _14849_/D vssd1 vssd1 vccd1 vccd1 _14849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08370_ hold711/A hold749/A hold579/A _14758_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08370_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_175_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07321_ _07332_/B _07321_/B _07321_/C vssd1 vssd1 vccd1 vccd1 _07321_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10256__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13602__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07252_ _08530_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08378_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2743_A _15177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07183_ hold2037/X _13651_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07183_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10019__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07903__A_N _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11508__C1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout403 _11643_/B vssd1 vssd1 vccd1 vccd1 _09925_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout414 _06978_/X vssd1 vssd1 vccd1 vccd1 _07010_/S sky130_fd_sc_hd__clkbuf_16
Xfanout425 _11877_/S vssd1 vssd1 vccd1 vccd1 _11893_/S sky130_fd_sc_hd__buf_8
XANTENNA_fanout394_A _07745_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _07710_/X vssd1 vssd1 vccd1 vccd1 _07742_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__08924__B1 _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__nand2_1
Xfanout447 _13792_/A2 vssd1 vssd1 vccd1 vccd1 _13625_/C sky130_fd_sc_hd__buf_4
Xfanout458 _12131_/X vssd1 vssd1 vccd1 vccd1 _12195_/A2 sky130_fd_sc_hd__buf_4
Xfanout469 _07884_/X vssd1 vssd1 vccd1 vccd1 _11640_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__07762__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ _09754_/B _09754_/C _09754_/A vssd1 vssd1 vccd1 vccd1 _09755_/Y sky130_fd_sc_hd__a21oi_1
X_06967_ _14083_/Q _06968_/C _06967_/C _14084_/Q vssd1 vssd1 vccd1 vccd1 _06967_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_119_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout561_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08706_ _08806_/B _08705_/C _08705_/A vssd1 vssd1 vccd1 vccd1 _08707_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09262__B _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09686_ _09547_/B _09549_/B _09683_/X _09685_/Y vssd1 vssd1 vccd1 vccd1 _09686_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_55_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _11645_/A _08637_/B vssd1 vssd1 vccd1 vccd1 _08637_/Y sky130_fd_sc_hd__nand2_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13028__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_A _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08568_ hold2732/X _12260_/A2 _12259_/A1 _13183_/B _08566_/Y vssd1 vssd1 vccd1 vccd1
+ _08568_/X sky130_fd_sc_hd__a221o_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12787__A1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07519_ hold2293/X _13690_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07519_/X sky130_fd_sc_hd__mux2_1
X_08499_ _08600_/B _08498_/C _08498_/A vssd1 vssd1 vccd1 vccd1 _08500_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ _10530_/A _10696_/B _10530_/C vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__nand3_2
XANTENNA__11313__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07002__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10463_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_49_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12200_ _12233_/A _12197_/X _12199_/X vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _13481_/A _13180_/B vssd1 vssd1 vccd1 vccd1 _15045_/D sky130_fd_sc_hd__and2_1
X_10392_ _10392_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12131_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12131_/X sky130_fd_sc_hd__or2_1
XFILLER_0_202_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12398__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__A2 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ _12128_/A hold2696/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12062_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07238__A _15226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold490 hold490/A vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08066__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _11011_/X _11013_/B vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12711__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07672__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ hold1837/X hold1621/X hold1599/X hold2301/X _12964_/S0 _13068_/A1 vssd1 vssd1
+ vccd1 vccd1 _12964_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08143__A1 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08143__B2 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 _11775_/X vssd1 vssd1 vccd1 vccd1 _14600_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12310__C _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _15377_/CLK hold912/X vssd1 vssd1 vccd1 vccd1 hold911/A sky130_fd_sc_hd__dfxtp_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _13703_/A1 hold1951/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A _12895_/B _13076_/A vssd1 vssd1 vccd1 vccd1 _12902_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_158_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11922__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _15369_/CLK _14634_/D vssd1 vssd1 vccd1 vccd1 _14634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ hold1431/X _15053_/Q _11861_/S vssd1 vssd1 vccd1 vccd1 _11846_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12778__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ hold697/X _13664_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 hold698/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14565_ _15435_/CLK hold220/X vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12873__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10728_ _10728_/A _10728_/B _10728_/C vssd1 vssd1 vccd1 vccd1 _10730_/A sky130_fd_sc_hd__or3_1
X_13516_ _13664_/A1 hold2295/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13516_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ _15264_/CLK hold940/X vssd1 vssd1 vccd1 vccd1 hold939/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _10836_/B _10658_/C _10658_/A vssd1 vssd1 vccd1 vccd1 _10660_/C sky130_fd_sc_hd__a21o_1
X_13447_ _09773_/B _13450_/A _13446_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15217_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12625__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11202__A1 _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11202__B2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ _13477_/A _13378_/B vssd1 vssd1 vccd1 vccd1 _15169_/D sky130_fd_sc_hd__and2_1
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08532__A _13384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ _15127_/CLK _15117_/D vssd1 vssd1 vccd1 vccd1 _15117_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10410__C1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12329_ _12329_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__and2_1
XANTENNA__10961__B1 _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12389__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15048_ _15369_/CLK _15048_/D vssd1 vssd1 vccd1 vccd1 _15048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2808 _14147_/Q vssd1 vssd1 vccd1 vccd1 hold2808/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_167_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12163__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2819 _15059_/Q vssd1 vssd1 vccd1 vccd1 hold2819/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13050__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _14091_/Q _06972_/C _07869_/X _06967_/X _06928_/Y vssd1 vssd1 vccd1 vccd1
+ _12301_/A sky130_fd_sc_hd__o32a_1
XFILLER_0_48_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07582__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09540_ _10129_/A _09708_/B _09429_/X _09430_/X _10142_/B vssd1 vssd1 vccd1 vccd1
+ _09545_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09471_ _09471_/A _09471_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _09471_/X sky130_fd_sc_hd__or3_1
XFILLER_0_176_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11832__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ _08317_/C _08318_/C _08519_/A _08421_/Y vssd1 vssd1 vccd1 vccd1 _08519_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_188_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13415__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__A1 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08353_ _13554_/A _08353_/B vssd1 vssd1 vccd1 vccd1 _08353_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12229__A _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07304_ _10022_/B _09858_/B vssd1 vssd1 vccd1 vccd1 _07305_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_132_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12864__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ _08269_/Y _08274_/Y _08283_/X _12241_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08285_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07235_ _08007_/A vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__inv_2
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout407_A _07149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07757__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07166_ _13519_/A0 hold2079/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07166_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07948__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ _13700_/A1 hold1549/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07097_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_A _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07492__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09807_ _13705_/A1 _11514_/A2 _11514_/B1 _13193_/B _09805_/Y vssd1 vssd1 vccd1 vccd1
+ _09807_/X sky130_fd_sc_hd__a221o_1
X_07999_ _08197_/A _07998_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _07999_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09738_ _09734_/Y _09735_/X _09590_/Y _09592_/X vssd1 vssd1 vccd1 vccd1 _09739_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_97_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ _10351_/A _10338_/C vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09873__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11742__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11700_ hold939/X _13654_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold940/A sky130_fd_sc_hd__mux2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _13080_/A1 _12679_/X _12677_/X vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__xnor2_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11562_ _11560_/X _11354_/B _11562_/S vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__mux2_1
X_14350_ _15378_/CLK hold408/X vssd1 vssd1 vccd1 vccd1 hold407/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13301_ input75/X fanout2/X _13300_/X vssd1 vssd1 vccd1 vccd1 _13302_/B sky130_fd_sc_hd__a21oi_1
X_10513_ _10513_/A _10513_/B _10513_/C vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__and3_1
XFILLER_0_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13669__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14281_ _15442_/CLK hold758/X vssd1 vssd1 vccd1 vccd1 hold757/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ _11493_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_190_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07667__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ hold553/X _13711_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold554/A sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__and2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13163_ _13390_/A _13163_/B vssd1 vssd1 vccd1 vccd1 _15028_/D sky130_fd_sc_hd__nor2_1
X_10375_ _10156_/X _10160_/B _10372_/Y _10374_/X vssd1 vssd1 vccd1 vccd1 _10439_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_21_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _12114_/A _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12114_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ _13100_/S0 _13089_/X _13093_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _13095_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12145__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ _12059_/A _12045_/B vssd1 vssd1 vccd1 vccd1 _14835_/D sky130_fd_sc_hd__and2_1
XANTENNA__11499__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09787__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13645__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13996_ _15394_/CLK _13996_/D vssd1 vssd1 vccd1 vccd1 _13996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ hold299/A hold431/A hold295/A _14742_/Q _12991_/S _13098_/S1 vssd1 vssd1
+ vccd1 vccd1 _12947_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_198_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _13673_/A1 _13103_/A2 _13078_/B1 _13194_/B vssd1 vssd1 vccd1 vccd1 _12878_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_160 _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13099__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07431__A _07431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_182 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13152__B _13152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_193 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ _15457_/CLK hold704/X vssd1 vssd1 vccd1 vccd1 hold703/A sky130_fd_sc_hd__dfxtp_1
X_11829_ _13716_/B _13683_/A vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12049__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12846__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14548_ _15452_/CLK _14548_/D vssd1 vssd1 vccd1 vccd1 _14548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09092__A2 _12275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14479_ _15062_/CLK _14479_/D vssd1 vssd1 vccd1 vccd1 _14479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07020_ hold2145/X _13691_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07020_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_141_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2441_A _15131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _09918_/A _13434_/B _08970_/X _10233_/A vssd1 vssd1 vccd1 vccd1 _08971_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13023__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2605 _14994_/Q vssd1 vssd1 vccd1 vccd1 hold2605/X sky130_fd_sc_hd__buf_2
XANTENNA__11827__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2616 _09093_/X vssd1 vssd1 vccd1 vccd1 _14439_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _13750_/A _13344_/B vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__nor2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2627 hold2830/X vssd1 vssd1 vccd1 vccd1 _10568_/B sky130_fd_sc_hd__clkbuf_2
Xhold2638 _12157_/X vssd1 vssd1 vccd1 vccd1 _14889_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1904 _11922_/X vssd1 vssd1 vccd1 vccd1 _14743_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2649 _14441_/Q vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1915 _14697_/Q vssd1 vssd1 vccd1 vccd1 hold1915/X sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ hold261/A _14066_/Q _14065_/Q hold573/A vssd1 vssd1 vccd1 vccd1 _07855_/C
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_78_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1926 _07625_/X vssd1 vssd1 vccd1 vccd1 _14248_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1937 _15268_/Q vssd1 vssd1 vccd1 vccd1 hold1937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1948 _13739_/X vssd1 vssd1 vccd1 vccd1 _15449_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1959 _14463_/Q vssd1 vssd1 vccd1 vccd1 hold1959/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07784_ hold1291/X _13689_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 _07784_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09523_ _09816_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _09533_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09821__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10967__A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13343__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09454_ _09454_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09454_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09950__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08405_ _09542_/A _08403_/X _08404_/X vssd1 vssd1 vccd1 vccd1 _08406_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ _10338_/B _09676_/D _09979_/C _10166_/A vssd1 vssd1 vccd1 vccd1 _09387_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout524_A _15425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08336_ _08380_/A _08333_/Y _08335_/C vssd1 vssd1 vccd1 vccd1 _08337_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12611__B1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08267_ _13870_/Q hold421/A hold905/A _13806_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08267_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_140_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07487__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07218_ _14056_/Q _14057_/Q hold573/A vssd1 vssd1 vccd1 vccd1 _07218_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ _14273_/Q hold801/A _14145_/Q _14463_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08199_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout893_A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08603__C _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07149_ _11928_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _07149_/X sky130_fd_sc_hd__or2_4
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10160_ _10160_/A _10160_/B _10160_/C vssd1 vssd1 vccd1 vccd1 _10336_/A sky130_fd_sc_hd__and3_1
XANTENNA__12127__C1 _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11737__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12678__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _14804_/Q hold649/A hold847/A _14740_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10092_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_22_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12773__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11350__B1 _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13850_ _15376_/CLK hold660/X vssd1 vssd1 vccd1 vccd1 hold659/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09153__D _15210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ _12951_/A _12801_/B vssd1 vssd1 vccd1 vccd1 _12802_/C sky130_fd_sc_hd__or2_1
XANTENNA__12525__S0 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _10992_/B _10992_/C _10992_/A vssd1 vssd1 vccd1 vccd1 _10994_/C sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_172_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13781_ hold163/X vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _13171_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _14957_/D sky130_fd_sc_hd__nor2_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07251__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15451_/CLK hold356/X vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12366_/A _12658_/X _12662_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12670_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _15435_/CLK hold410/X vssd1 vssd1 vccd1 vccd1 hold409/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07609__A0 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _11614_/A _11614_/B vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11204__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_187_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ _15382_/CLK hold844/X vssd1 vssd1 vccd1 vccd1 hold843/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12700_/S0 _12589_/X _12593_/X _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12595_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ _15434_/CLK hold596/X vssd1 vssd1 vccd1 vccd1 hold595/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11545_ _11545_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11546_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08282__B1 _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15408_/CLK sky130_fd_sc_hd__clkbuf_16
X_11476_ _13749_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _11476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14264_ _15068_/CLK _14264_/D vssd1 vssd1 vccd1 vccd1 _14264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_110_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12905__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ _14678_/Q _13951_/Q hold437/A _13919_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10428_/B sky130_fd_sc_hd__mux4_1
X_13215_ hold1031/X _13727_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13215_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09231__C1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14195_ _15190_/CLK hold168/X vssd1 vssd1 vccd1 vccd1 _14195_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10916__B1 _10951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09782__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _10700_/A _11542_/B _10524_/A _10358_/D vssd1 vssd1 vccd1 vccd1 _10524_/B
+ sky130_fd_sc_hd__nand4_2
X_13146_ _13381_/A _13146_/B vssd1 vssd1 vccd1 vccd1 _15011_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08810__A _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13102_/A _13077_/B _13077_/C vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__and3_1
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__xor2_2
XANTENNA_clkbuf_leaf_125_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13330__A1 input150/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12028_ hold2562/X hold2718/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12028_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12764__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__B _13147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11892__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09641__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13979_ _15379_/CLK _13979_/D vssd1 vssd1 vccd1 vccd1 _13979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__D _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07943__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__A2_N _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ _10183_/A _09979_/B _09712_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _09297_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08121_ _08197_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_122_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08052_ _13867_/Q hold387/A _13835_/Q _13803_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08052_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_141_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07100__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ _13675_/A1 hold1481/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07003_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09816__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__D _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13338__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2402 hold2839/X vssd1 vssd1 vccd1 vccd1 _08179_/B sky130_fd_sc_hd__buf_1
Xinput109 in1[20] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__clkbuf_1
X_08954_ _08997_/B _08954_/B _08955_/B vssd1 vssd1 vccd1 vccd1 _08954_/X sky130_fd_sc_hd__and3_1
Xhold2413 _15036_/Q vssd1 vssd1 vccd1 vccd1 _07576_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2424 _14856_/Q vssd1 vssd1 vccd1 vccd1 hold2424/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13321__A1 input147/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__B1 _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2435 _14853_/Q vssd1 vssd1 vccd1 vccd1 hold2435/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ _07904_/A _07904_/B _07430_/A vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__a21o_1
Xhold2446 _15459_/Q vssd1 vssd1 vccd1 vccd1 _13536_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1701 _13839_/Q vssd1 vssd1 vccd1 vccd1 hold1701/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1712 _07122_/X vssd1 vssd1 vccd1 vccd1 _13932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2457 _14855_/Q vssd1 vssd1 vccd1 vccd1 hold2457/X sky130_fd_sc_hd__dlygate4sd3_1
X_08885_ _09164_/A _09860_/B _08804_/A _08801_/X vssd1 vssd1 vccd1 vccd1 _08950_/A
+ sky130_fd_sc_hd__a31o_1
Xhold2468 _12113_/X vssd1 vssd1 vccd1 vccd1 _14868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1723 _13879_/Q vssd1 vssd1 vccd1 vccd1 hold1723/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11332__B1 _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1734 _07120_/X vssd1 vssd1 vccd1 vccd1 _13930_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2479 _09926_/X vssd1 vssd1 vccd1 vccd1 _14445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 _13877_/Q vssd1 vssd1 vccd1 vccd1 hold1745/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1756 _11876_/X vssd1 vssd1 vccd1 vccd1 _14698_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07836_ _07819_/X _07826_/Y _07835_/X _12241_/A vssd1 vssd1 vccd1 vccd1 _07882_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1767 _15390_/Q vssd1 vssd1 vccd1 vccd1 hold1767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1778 _11674_/X vssd1 vssd1 vccd1 vccd1 _14477_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07770__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1789 _13878_/Q vssd1 vssd1 vccd1 vccd1 hold1789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout641_A _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _13738_/A1 hold1963/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07767_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13624__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout739_A _14954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08187__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09506_ _09941_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__or2_1
XANTENNA__10438__A2 _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07698_ hold1871/X _13671_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09701__D _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09437_/A _09712_/B _09437_/C _09437_/D vssd1 vssd1 vccd1 vccd1 _09437_/Y
+ sky130_fd_sc_hd__nand4_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _10244_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08319_ _08318_/B _08318_/C _08318_/A vssd1 vssd1 vccd1 vccd1 _08320_/D sky130_fd_sc_hd__a21oi_1
X_09299_ _09979_/B _10022_/B _09858_/C _09542_/A vssd1 vssd1 vccd1 vccd1 _09301_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11494__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15411_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_60 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11330_ _11330_/A vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__inv_2
XFILLER_0_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_82 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_93 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10610__A2 _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07010__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11040__B _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _11329_/B _11259_/X _11029_/X _11033_/C vssd1 vssd1 vccd1 vccd1 _11261_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08567__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ _10058_/Y _10060_/Y _10386_/B _10211_/X vssd1 vssd1 vccd1 vccd1 _10392_/A
+ sky130_fd_sc_hd__a211oi_2
X_13000_ _12996_/X _12997_/X _12999_/X _12998_/X _13050_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _13001_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09726__A _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _11192_/A _11192_/B vssd1 vssd1 vccd1 vccd1 _11200_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_63_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13248__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ _10142_/B _14956_/Q _14957_/Q _11573_/A vssd1 vssd1 vccd1 vccd1 _10144_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09445__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__A1 input144/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12115__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12746__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _10265_/A _10073_/C _10073_/A vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__a21oi_1
X_14951_ _15222_/CLK _14951_/D vssd1 vssd1 vccd1 vccd1 _14951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13682__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ _15435_/CLK _13902_/D vssd1 vssd1 vccd1 vccd1 _13902_/Q sky130_fd_sc_hd__dfxtp_1
X_14882_ _14889_/CLK _14882_/D vssd1 vssd1 vccd1 vccd1 _14882_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07680__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _15072_/CLK _13833_/D vssd1 vssd1 vccd1 vccd1 _13833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ hold219/X vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__clkbuf_1
X_10976_ _10976_/A _10976_/B _10791_/Y vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__or3b_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ _14410_/Q _14122_/Q _12741_/S vssd1 vssd1 vccd1 vccd1 _12715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ hold777/X _13728_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 hold778/A sky130_fd_sc_hd__mux2_1
XANTENNA__11930__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15434_ _15434_/CLK _15434_/D vssd1 vssd1 vccd1 vccd1 _15434_/Q sky130_fd_sc_hd__dfxtp_1
X_12646_ hold459/A _15274_/Q hold927/A _14375_/Q _12641_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12646_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_183_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13430__B _13430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15365_ _15365_/CLK hold648/X vssd1 vssd1 vccd1 vccd1 hold647/A sky130_fd_sc_hd__dfxtp_1
X_12577_ _13027_/A _12577_/B _12577_/C vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__and3_1
XANTENNA__12327__A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14316_ _15410_/CLK _14316_/D vssd1 vssd1 vccd1 vccd1 _14316_/Q sky130_fd_sc_hd__dfxtp_1
X_11528_ _11528_/A _11528_/B vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ _15296_/CLK _15296_/D vssd1 vssd1 vccd1 vccd1 _15296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 hold319/A vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14247_ _15405_/CLK _14247_/D vssd1 vssd1 vccd1 vccd1 _14247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _11459_/A _11459_/B vssd1 vssd1 vccd1 vccd1 _11461_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14178_ _15179_/CLK hold152/X vssd1 vssd1 vccd1 vccd1 _14178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08653__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13129_/A hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__and2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13303__A1 input141/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _07504_/X vssd1 vssd1 vccd1 vccd1 _14132_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1019 _13828_/Q vssd1 vssd1 vccd1 vccd1 hold1019/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08670_ _08776_/B _09860_/A vssd1 vssd1 vccd1 vccd1 _08674_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07590__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07621_ hold831/X _13727_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 hold832/A sky130_fd_sc_hd__mux2_1
XANTENNA__13067__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07552_ _13393_/A hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__and2_1
XFILLER_0_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08494__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07483_ hold1113/X _13689_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07483_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _09350_/B _09222_/B vssd1 vssd1 vccd1 vccd1 _09222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09153_ _10166_/A _11333_/B _09709_/B _15210_/Q vssd1 vssd1 vccd1 vccd1 _09154_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__08246__B1 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11141__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08104_ _07900_/B _13379_/B _08072_/X vssd1 vssd1 vccd1 vccd1 _13416_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_185_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _09082_/X _09084_/B vssd1 vssd1 vccd1 vccd1 _09086_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08035_ _07976_/A _07975_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_142_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput80 in0[23] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_1
XANTENNA__10980__A _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 hold820/A vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput91 in0[4] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_1
XFILLER_0_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08549__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 hold831/A vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07765__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 hold842/A vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 hold853/A vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold864 hold864/A vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 hold875/A vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11287__S _11287_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 hold886/A vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold897 hold897/A vssd1 vssd1 vccd1 vccd1 hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _09987_/A _09987_/B _09987_/C vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__and3_1
XFILLER_0_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2210 _07086_/X vssd1 vssd1 vccd1 vccd1 _13899_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2221 _14030_/Q vssd1 vssd1 vccd1 vccd1 _07455_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2232 _07130_/X vssd1 vssd1 vccd1 vccd1 _13940_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ _08817_/Y _08819_/X _08935_/X _08936_/Y vssd1 vssd1 vccd1 vccd1 _08940_/B
+ sky130_fd_sc_hd__o211ai_4
Xhold2243 _14382_/Q vssd1 vssd1 vccd1 vccd1 hold2243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06980__A0 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2254 _11929_/X vssd1 vssd1 vccd1 vccd1 _14749_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1520 _13663_/X vssd1 vssd1 vccd1 vccd1 _15370_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2265 _14537_/Q vssd1 vssd1 vccd1 vccd1 hold2265/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1531 _14112_/Q vssd1 vssd1 vccd1 vccd1 hold1531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2276 _13472_/X vssd1 vssd1 vccd1 vccd1 _15231_/D sky130_fd_sc_hd__buf_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1542 _13219_/X vssd1 vssd1 vccd1 vccd1 _15083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2287 _13902_/Q vssd1 vssd1 vccd1 vccd1 hold2287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ hold639/A _14507_/Q hold887/A _14731_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08869_/B sky130_fd_sc_hd__mux4_1
Xhold1553 _14349_/Q vssd1 vssd1 vccd1 vccd1 hold1553/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2298 _07072_/X vssd1 vssd1 vccd1 vccd1 _13888_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 _07085_/X vssd1 vssd1 vccd1 vccd1 _13898_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09281__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1575 _14785_/Q vssd1 vssd1 vccd1 vccd1 hold1575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1586 _11905_/X vssd1 vssd1 vccd1 vccd1 _14726_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07819_ _12243_/A _07815_/Y _07817_/Y _07818_/Y vssd1 vssd1 vccd1 vccd1 _07819_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1597 _14229_/Q vssd1 vssd1 vccd1 vccd1 hold1597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08799_ _08799_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08800_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10830_ _14952_/Q _10830_/B _10830_/C _10830_/D vssd1 vssd1 vccd1 vccd1 _10830_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07005__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12900__S0 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _15385_/Q _15288_/Q hold553/A _14389_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10761_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11750__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _12496_/X _12497_/X _12499_/X _12498_/X _12644_/A1 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12501_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_165_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ _11567_/A _15223_/Q vssd1 vssd1 vccd1 vccd1 _10694_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10831__A2 _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13480_ _13492_/A hold123/X vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__and2_1
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12569__C1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _08038_/B _08636_/A _13144_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12432_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15150_ _15313_/CLK _15150_/D vssd1 vssd1 vccd1 vccd1 _15150_/Q sky130_fd_sc_hd__dfxtp_1
X_12362_ hold453/A hold975/A hold635/A _13896_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12362_/X sky130_fd_sc_hd__mux4_1
X_14101_ _14105_/CLK hold258/X vssd1 vssd1 vccd1 vccd1 _14101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13677__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10595__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _11497_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/Y sky130_fd_sc_hd__nor2_1
X_12293_ _15347_/Q _15346_/Q vssd1 vssd1 vccd1 vccd1 _13240_/C sky130_fd_sc_hd__nor2_1
X_15081_ _15440_/CLK _15081_/D vssd1 vssd1 vccd1 vccd1 _15081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07675__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ _11351_/B _11586_/B _11620_/B _11541_/A vssd1 vssd1 vccd1 vccd1 _11247_/C
+ sky130_fd_sc_hd__a22o_1
X_14032_ _15293_/CLK _14032_/D vssd1 vssd1 vccd1 vccd1 _14032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11544__B1 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07212__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ _10987_/D _10987_/Y _11173_/Y _11174_/X vssd1 vssd1 vccd1 vccd1 _11177_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _10126_/A _10126_/B _11606_/A vssd1 vssd1 vccd1 vccd1 _10126_/X sky130_fd_sc_hd__and3_1
XFILLER_0_98_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output239_A _15460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _10056_/A _10056_/B _10056_/C _10056_/D vssd1 vssd1 vccd1 vccd1 _10057_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14934_ _15256_/CLK _14934_/D vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14865_ _14866_/CLK _14865_/D vssd1 vssd1 vccd1 vccd1 _14865_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13816_ _15087_/CLK _13816_/D vssd1 vssd1 vccd1 vccd1 _13816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14796_ _15373_/CLK hold938/X vssd1 vssd1 vccd1 vccd1 hold937/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13747_ hold399/X hold2817/X _13748_/S vssd1 vssd1 vccd1 vccd1 hold400/A sky130_fd_sc_hd__mux2_1
X_10959_ _10268_/A _10268_/B _10736_/Y _10958_/X vssd1 vssd1 vccd1 vccd1 _10959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11660__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13441__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08535__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13678_ hold1365/X _15064_/Q _13682_/S vssd1 vssd1 vccd1 vccd1 _13678_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10784__B _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13160__B _13160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15417_ _15454_/CLK _15417_/D vssd1 vssd1 vccd1 vccd1 _15417_/Q sky130_fd_sc_hd__dfxtp_1
X_12629_ _13386_/B _12325_/B _12628_/X vssd1 vssd1 vccd1 vccd1 _12629_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__A1 _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__B2 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15348_ _15348_/CLK _15348_/D vssd1 vssd1 vccd1 vccd1 _15348_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08874__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__S _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15376_/CLK _15279_/D vssd1 vssd1 vccd1 vccd1 _15279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07585__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10008__C _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09366__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12958__S0 _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ _09839_/B _09839_/C _09839_/A vssd1 vssd1 vccd1 vccd1 _09841_/C sky130_fd_sc_hd__o21ai_1
Xfanout607 _11407_/A vssd1 vssd1 vccd1 vccd1 _11605_/A sky130_fd_sc_hd__clkbuf_8
Xfanout618 _15205_/Q vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2619_A _14431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout629 _15202_/Q vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10305__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _11288_/A1 _13394_/B _09654_/X vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__a21oi_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _13655_/A1 hold929/X _06994_/S vssd1 vssd1 vccd1 vccd1 hold930/A sky130_fd_sc_hd__mux2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11835__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ _08721_/B _08721_/C _08680_/X vssd1 vssd1 vccd1 vccd1 _08722_/X sky130_fd_sc_hd__a21bo_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _14793_/Q _14505_/Q _14633_/Q _14729_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08654_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10678__C _15219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07604_ _13743_/A1 hold1621/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07604_/X sky130_fd_sc_hd__mux2_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08584_ _09026_/B _09437_/A _08685_/C _08908_/A vssd1 vssd1 vccd1 vccd1 _08586_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07535_ hold691/X hold2819/X _07544_/S vssd1 vssd1 vccd1 vccd1 hold692/A sky130_fd_sc_hd__mux2_1
XANTENNA__08467__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12666__S _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout437_A _07644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ _13501_/A hold37/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__and2_1
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09205_ _09205_/A _09205_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09205_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07397_ hold255/X _07450_/B vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__and2_1
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout604_A _15209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _09136_/A _09253_/A _09714_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09138_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _08916_/X _08919_/X _09065_/A _09066_/X vssd1 vssd1 vccd1 vccd1 _09199_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_161_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07495__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ _08091_/A _08017_/B _08017_/C vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12949__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold650 hold650/A vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 hold661/A vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 hold672/A vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10860__D _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold683 hold683/A vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 hold694/A vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ _14942_/Q _10338_/C _09817_/A _09814_/X vssd1 vssd1 vccd1 vccd1 _09971_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2040 _07652_/X vssd1 vssd1 vccd1 vccd1 _14273_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2051 _14378_/Q vssd1 vssd1 vccd1 vccd1 hold2051/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11745__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2062 _11918_/X vssd1 vssd1 vccd1 vccd1 _14739_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2073 _15286_/Q vssd1 vssd1 vccd1 vccd1 hold2073/X sky130_fd_sc_hd__dlygate4sd3_1
X_12980_ _13080_/A1 _12979_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _12980_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2084 _07135_/X vssd1 vssd1 vccd1 vccd1 _13945_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__B _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2095 _13906_/Q vssd1 vssd1 vccd1 vccd1 hold2095/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1350 _07074_/X vssd1 vssd1 vccd1 vccd1 _13890_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1361 _13970_/Q vssd1 vssd1 vccd1 vccd1 hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1372 _07760_/X vssd1 vssd1 vccd1 vccd1 _14376_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ _13719_/A1 hold1179/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 _14637_/Q vssd1 vssd1 vccd1 vccd1 hold1383/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _11683_/X vssd1 vssd1 vccd1 vccd1 _14486_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _15387_/CLK hold728/X vssd1 vssd1 vccd1 vccd1 hold727/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11862_ _13716_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _11894_/S sky130_fd_sc_hd__nor2_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13601_ input44/X _13634_/B _13625_/B vssd1 vssd1 vccd1 vccd1 _15327_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_184_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11057__A2 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10813_ _10978_/B _10812_/C _10812_/A vssd1 vssd1 vccd1 vccd1 _10814_/C sky130_fd_sc_hd__a21o_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14581_ _14581_/CLK hold280/X vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__dfxtp_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ hold1033/X _13746_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_200_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ _13680_/A1 hold1145/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ _10744_/A _10744_/B vssd1 vssd1 vccd1 vccd1 _10745_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_211_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _13535_/B _13463_/B vssd1 vssd1 vccd1 vccd1 _15225_/D sky130_fd_sc_hd__and2_1
X_10675_ _10502_/B _10502_/Y _10673_/Y _10674_/X vssd1 vssd1 vccd1 vccd1 _10675_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08074__B _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ _15324_/CLK hold444/X vssd1 vssd1 vccd1 vccd1 _15202_/Q sky130_fd_sc_hd__dfxtp_4
X_12414_ _14270_/Q _14206_/Q hold751/A hold1631/X _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12414_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13754__A1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13394_ _13397_/A _13394_/B vssd1 vssd1 vccd1 vccd1 _15185_/D sky130_fd_sc_hd__and2_1
XFILLER_0_211_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output189_A _15170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _15460_/CLK _15133_/D vssd1 vssd1 vccd1 vccd1 _15133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12345_ _12692_/A1 _12344_/X _12343_/X _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12345_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12309__A2 _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15064_ _15196_/CLK _15064_/D vssd1 vssd1 vccd1 vccd1 _15064_/Q sky130_fd_sc_hd__dfxtp_1
X_12276_ _13389_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _14925_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _15382_/CLK _14015_/D vssd1 vssd1 vccd1 vccd1 _14015_/Q sky130_fd_sc_hd__dfxtp_1
X_11227_ _11224_/Y _11337_/A _11335_/A _15224_/Q vssd1 vssd1 vccd1 vccd1 _11337_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_103_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__B _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _11158_/A _11158_/B _11158_/C vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_65_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11655__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10109_ _10002_/C _10108_/C _14963_/Q _11578_/A vssd1 vssd1 vccd1 vccd1 _10110_/D
+ sky130_fd_sc_hd__a22o_1
X_11089_ _11089_/A _11089_/B _11089_/C vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__or3_1
XFILLER_0_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13155__B _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ _14926_/CLK _14917_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12493__A1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _14975_/CLK _14848_/D vssd1 vssd1 vccd1 vccd1 _14848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14779_ _15287_/CLK hold796/X vssd1 vssd1 vccd1 vccd1 hold795/A sky130_fd_sc_hd__dfxtp_1
X_07320_ _09767_/A _07320_/B _09914_/B _07320_/D vssd1 vssd1 vccd1 vccd1 _07321_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_128_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12340__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ _09712_/A _09858_/A vssd1 vssd1 vccd1 vccd1 _08527_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold2471_A _14989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07672__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07182_ _07182_/A _11730_/A vssd1 vssd1 vccd1 vccd1 _07182_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11756__A0 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10019__B _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout404 _11643_/B vssd1 vssd1 vccd1 vccd1 _07812_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__10035__A _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 _13716_/Y vssd1 vssd1 vccd1 vccd1 _13732_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout426 _11894_/S vssd1 vssd1 vccd1 vccd1 _11877_/S sky130_fd_sc_hd__buf_12
XANTENNA__08924__B2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _09720_/A _09719_/B _09717_/X vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__a21o_1
Xfanout437 _07644_/Y vssd1 vssd1 vccd1 vccd1 _07660_/S sky130_fd_sc_hd__buf_12
Xfanout448 _07389_/Y vssd1 vssd1 vccd1 vccd1 _13792_/A2 sky130_fd_sc_hd__buf_4
Xfanout459 _12194_/B vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout387_A _11696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13346__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _09754_/A _09754_/B _09754_/C vssd1 vssd1 vccd1 vccd1 _09754_/X sky130_fd_sc_hd__and3_1
XANTENNA__09543__B _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06966_ _14081_/Q _14085_/Q vssd1 vssd1 vccd1 vccd1 _06967_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08705_ _08705_/A _08806_/B _08705_/C vssd1 vssd1 vccd1 vccd1 _08805_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09262__C _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ _09684_/B _09684_/C _09684_/A vssd1 vssd1 vccd1 vccd1 _09685_/Y sky130_fd_sc_hd__a21oi_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_A _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15254_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _08636_/A vssd1 vssd1 vccd1 vccd1 _08636_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_179_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10590__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout721_A _14964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ hold2753/X input3/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13183_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_A _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ hold1679/X _13689_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07518_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08498_ _08498_/A _08600_/B _08498_/C vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08175__A _13380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07449_ hold127/X _07450_/B vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__and2_1
XFILLER_0_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12128__C _12128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ _10460_/A _10460_/B vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12944__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _09119_/A _09119_/B _09119_/C vssd1 vssd1 vccd1 vccd1 _09119_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_126_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10391_ _10560_/B _10391_/B vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__or2_1
XFILLER_0_150_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09168__B2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _12063_/A _12061_/B vssd1 vssd1 vccd1 vccd1 _14843_/D sky130_fd_sc_hd__and2_1
XANTENNA__07238__B _14970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12398__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07179__A0 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 hold480/A vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 hold491/A vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ _11008_/X _11010_/Y _10826_/X _10829_/X vssd1 vssd1 vccd1 vccd1 _11013_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07254__A _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ _06943_/A _12958_/X _12962_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12970_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13690__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15385_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1180 _11931_/X vssd1 vssd1 vccd1 vccd1 _14751_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08143__A2 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _15439_/CLK _14702_/D vssd1 vssd1 vccd1 vccd1 _14702_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1191 _14599_/Q vssd1 vssd1 vccd1 vccd1 hold1191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__B1 _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ _13669_/A1 hold2047/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _13050_/S0 _12889_/X _12893_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _12895_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _15440_/CLK _14633_/D vssd1 vssd1 vccd1 vccd1 _14633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ hold1247/X _13732_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12778__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11504__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14564_ _15264_/CLK hold180/X vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__dfxtp_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ hold1195/X _13663_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11776_/X sky130_fd_sc_hd__mux2_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13515_ _13663_/A1 hold1845/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__mux2_1
X_10727_ _10723_/Y _10724_/X _10553_/B _10552_/Y vssd1 vssd1 vccd1 vccd1 _10728_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14495_ _15263_/CLK _14495_/D vssd1 vssd1 vccd1 vccd1 _14495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13446_ _13450_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _13446_/Y sky130_fd_sc_hd__nand2_1
X_10658_ _10658_/A _10836_/B _10658_/C vssd1 vssd1 vccd1 vccd1 _10660_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11738__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11202__A2 _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13377_ _13477_/A _13377_/B vssd1 vssd1 vccd1 vccd1 _15168_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10589_ _11497_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10589_/Y sky130_fd_sc_hd__nor2_1
X_15116_ _15116_/CLK _15116_/D vssd1 vssd1 vccd1 vccd1 _15116_/Q sky130_fd_sc_hd__dfxtp_1
X_12328_ _12601_/A _12316_/Y _12322_/Y _12327_/A vssd1 vssd1 vccd1 vccd1 _12328_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10961__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__B2 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ _15079_/CLK _15047_/D vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__dfxtp_1
X_12259_ _12259_/A1 _13173_/B _13375_/B _07900_/B vssd1 vssd1 vccd1 vccd1 _12259_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2809 _15065_/Q vssd1 vssd1 vccd1 vccd1 hold2809/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13166__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15418_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_204_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08765__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09470_ _09471_/A _09471_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _09470_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_188_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08421_ _08516_/A _08420_/C _08420_/A vssd1 vssd1 vccd1 vccd1 _08421_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13613__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11414__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08352_ _13554_/A _08352_/B _08352_/C vssd1 vssd1 vccd1 vccd1 _08544_/C sky130_fd_sc_hd__and3_1
XFILLER_0_59_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12313__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07103__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07303_ _10022_/B _09858_/B vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__and2_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12520__C_N _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ _08880_/A1 _08276_/Y _08278_/Y _08280_/Y _08282_/Y vssd1 vssd1 vccd1 vccd1
+ _08283_/X sky130_fd_sc_hd__o32a_1
X_07234_ _08075_/B _11566_/A vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07165_ _13666_/A1 hold1319/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07165_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12245__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12670__C_N _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _13732_/A1 hold1681/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07096_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07773__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout769_A _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ hold2763/X input14/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__mux2_2
XANTENNA__13076__A _13076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07581__A0 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ _15394_/Q _14529_/Q hold671/A _14753_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07998_/X sky130_fd_sc_hd__mux4_1
X_09737_ _09590_/Y _09592_/X _09734_/Y _09735_/X vssd1 vssd1 vccd1 vccd1 _09739_/B
+ sky130_fd_sc_hd__a211o_1
X_06949_ _14036_/Q hold273/A hold237/A vssd1 vssd1 vccd1 vccd1 _06950_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_66_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _15229_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08756__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08619_ _08508_/Y _08510_/Y _08617_/Y _08618_/X vssd1 vssd1 vccd1 vccd1 _08621_/B
+ sky130_fd_sc_hd__a211oi_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09599_ _09599_/A _09599_/B _09599_/C vssd1 vssd1 vccd1 vccd1 _09601_/C sky130_fd_sc_hd__or3_4
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13015__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11630_ _11630_/A _11630_/B vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__xnor2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07013__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11561_ _11561_/A _15221_/Q vssd1 vssd1 vccd1 vccd1 _11562_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ input139/X fanout5/X fanout3/X input107/X vssd1 vssd1 vccd1 vccd1 _13300_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13709__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ _11335_/A _11586_/B _10340_/B _10338_/X vssd1 vssd1 vccd1 vccd1 _10513_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07948__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14280_ _14791_/CLK hold800/X vssd1 vssd1 vccd1 vccd1 hold799/A sky130_fd_sc_hd__dfxtp_1
X_11492_ _14361_/Q _14265_/Q hold885/A _14137_/Q _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _11493_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_162_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13231_ hold523/X hold2765/A _13236_/S vssd1 vssd1 vccd1 vccd1 hold524/A sky130_fd_sc_hd__mux2_1
X_10443_ _10443_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13162_ _13390_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _15027_/D sky130_fd_sc_hd__nor2_1
X_10374_ _10373_/B _10373_/C _10373_/A vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13685__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ hold2467/X _12129_/A2 _12112_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12113_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ _13098_/S1 _13090_/X _13092_/X vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07683__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ hold2553/X hold2705/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout790 _12601_/A vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13995_ _14754_/CLK hold388/X vssd1 vssd1 vccd1 vccd1 hold387/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_57_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15116_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11933__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _15383_/Q _15286_/Q hold393/A _14387_/Q _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12946_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_88_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_150 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _13102_/A _12877_/B _12877_/C vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__and3_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_161 _15423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_172 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14616_ _15385_/CLK hold624/X vssd1 vssd1 vccd1 vccd1 hold623/A sky130_fd_sc_hd__dfxtp_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_183 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ hold787/X _13715_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold788/A sky130_fd_sc_hd__mux2_1
XFILLER_0_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_194 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _15449_/CLK _14547_/D vssd1 vssd1 vccd1 vccd1 _14547_/Q sky130_fd_sc_hd__dfxtp_1
X_11759_ _13745_/A1 hold1491/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09639__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14478_ _15063_/CLK hold730/X vssd1 vssd1 vccd1 vccd1 hold729/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13429_ _08640_/A _13440_/S _13428_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _13429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08970_ _15147_/Q _09925_/A2 _08256_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _08970_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07593__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2606 _12175_/X vssd1 vssd1 vccd1 vccd1 _14898_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07921_ _07921_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12687__A1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2617 _14983_/Q vssd1 vssd1 vccd1 vccd1 hold2617/X sky130_fd_sc_hd__buf_2
XFILLER_0_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2628 _14977_/Q vssd1 vssd1 vccd1 vccd1 hold2628/X sky130_fd_sc_hd__buf_2
Xhold2639 _15138_/Q vssd1 vssd1 vccd1 vccd1 hold2639/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08986__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1905 _14220_/Q vssd1 vssd1 vccd1 vccd1 hold1905/X sky130_fd_sc_hd__dlygate4sd3_1
X_07852_ _07852_/A _07852_/B vssd1 vssd1 vccd1 vccd1 _07857_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12004__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1916 _11875_/X vssd1 vssd1 vccd1 vccd1 _14697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1927 _14480_/Q vssd1 vssd1 vccd1 vccd1 hold1927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1938 _13510_/X vssd1 vssd1 vccd1 vccd1 _15268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1949 _14595_/Q vssd1 vssd1 vccd1 vccd1 hold1949/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput1 dmemresp_rdata[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_07783_ hold779/X _13721_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold780/A sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15348_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11843__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _09393_/A _09392_/B _09392_/A vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_127_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09821__B _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__B _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _09454_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09453_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08404_ _08776_/A _08809_/B _08809_/D _09008_/A vssd1 vssd1 vccd1 vccd1 _08404_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11144__A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09384_ _09661_/A _09979_/D vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08335_ _08380_/A _08335_/B _08335_/C vssd1 vssd1 vccd1 vccd1 _08380_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12611__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout517_A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10622__B1 _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ hold219/A _14306_/Q _14597_/Q _13966_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08266_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07217_ hold255/X hold271/A hold313/A hold281/A vssd1 vssd1 vccd1 vccd1 _07855_/A
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08197_ _08197_/A _08197_/B vssd1 vssd1 vccd1 vccd1 _08197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08603__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ _14088_/Q _14089_/Q _14090_/Q vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__or3_4
XFILLER_0_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07079_ _07744_/A _11729_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__or3_2
XFILLER_0_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09284__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ _15381_/Q _15284_/Q _15092_/Q _14385_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10090_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12678__B2 _13186_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12773__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A1 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__B2 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07008__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _14954_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11753__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _12796_/X _12797_/X _12799_/X _12798_/X _12844_/A1 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12801_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12525__S1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ hold279/X vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11102__A1 _06941_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ _10992_/A _10992_/B _10992_/C vssd1 vssd1 vccd1 vccd1 _10994_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _13106_/A1 _13156_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__o21a_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11054__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__B1 _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15450_ _15450_/CLK hold330/X vssd1 vssd1 vccd1 vccd1 hold329/A sky130_fd_sc_hd__dfxtp_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12662_ _12668_/A1 _12659_/X _12661_/X vssd1 vssd1 vccd1 vccd1 _12662_/X sky130_fd_sc_hd__a21o_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14401_ _15040_/CLK hold442/X vssd1 vssd1 vccd1 vccd1 hold441/A sky130_fd_sc_hd__dfxtp_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11613_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__xnor2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12584__S _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ _15408_/CLK _15381_/D vssd1 vssd1 vccd1 vccd1 _15381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ _12699_/S1 _12590_/X _12592_/X vssd1 vssd1 vccd1 vccd1 _12593_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11204__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07678__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14332_ _15392_/CLK hold526/X vssd1 vssd1 vccd1 vccd1 hold525/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08282__A1 _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ _11420_/X _11449_/A _11390_/A _11378_/C vssd1 vssd1 vccd1 vccd1 _11545_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08363__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14263_ _14909_/CLK hold798/X vssd1 vssd1 vccd1 vccd1 hold797/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11475_ _07879_/X _13404_/B _11322_/X vssd1 vssd1 vccd1 vccd1 _13466_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_162_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13563__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ hold889/X _13512_/A0 _13220_/S vssd1 vssd1 vccd1 vccd1 hold890/A sky130_fd_sc_hd__mux2_1
XFILLER_0_123_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10426_ _10426_/A _10426_/B vssd1 vssd1 vccd1 vccd1 _10426_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14194_ _15190_/CLK hold162/X vssd1 vssd1 vccd1 vccd1 _14194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output171_A _15183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _13381_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _15010_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10357_ _11351_/B _10356_/C _11536_/B _14947_/Q vssd1 vssd1 vccd1 vccd1 _10358_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08810__B _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13428__B _13428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12669__A1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12213__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ _13076_/A _13076_/B vssd1 vssd1 vccd1 vccd1 _13077_/C sky130_fd_sc_hd__or2_1
X_10288_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10463_/B sky130_fd_sc_hd__nor2_1
X_12027_ _12063_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _14826_/D sky130_fd_sc_hd__and2_1
XFILLER_0_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12764__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09922__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12759__S _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13094__A1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ _15376_/CLK _13978_/D vssd1 vssd1 vccd1 vccd1 _13978_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07442__A _08107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__B _13163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ _13398_/B _13104_/A2 _12928_/X vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_76_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08257__B _14430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07943__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07588__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08120_ _14787_/Q _14499_/Q hold995/A _14723_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08121_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10080__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ hold263/A _14303_/Q _14594_/Q _13963_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08051_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07002_ _13674_/A1 hold867/X _07010_/S vssd1 vssd1 vccd1 vccd1 hold868/A sky130_fd_sc_hd__mux2_1
XFILLER_0_4_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08120__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__B _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08953_ _08953_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08955_/B sky130_fd_sc_hd__or2_1
XFILLER_0_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2403 _13549_/X vssd1 vssd1 vccd1 vccd1 _15300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2414 _14059_/Q vssd1 vssd1 vccd1 vccd1 _06918_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09525__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2425 _12089_/X vssd1 vssd1 vccd1 vccd1 _14856_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07904_ _07904_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _08036_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2436 _12083_/X vssd1 vssd1 vccd1 vccd1 _14853_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09525__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1702 _07022_/X vssd1 vssd1 vccd1 vccd1 _13839_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2447 _15340_/Q vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08884_ _13698_/A1 _11514_/A2 _11514_/B1 _13186_/B _08882_/Y vssd1 vssd1 vccd1 vccd1
+ _08884_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11332__A1 _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1713 _14368_/Q vssd1 vssd1 vccd1 vccd1 hold1713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2458 _12087_/X vssd1 vssd1 vccd1 vccd1 _14855_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11332__B2 _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1724 _07063_/X vssd1 vssd1 vccd1 vccd1 _13879_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10766__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2469 _14854_/Q vssd1 vssd1 vccd1 vccd1 hold2469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1735 _14400_/Q vssd1 vssd1 vccd1 vccd1 hold1735/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07835_ _06926_/A _07828_/Y _07830_/Y _07832_/Y _07834_/Y vssd1 vssd1 vccd1 vccd1
+ _07835_/X sky130_fd_sc_hd__o32a_1
Xhold1746 _07061_/X vssd1 vssd1 vccd1 vccd1 _13877_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1757 _15092_/Q vssd1 vssd1 vccd1 vccd1 hold1757/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout467_A _11287_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1768 _13684_/X vssd1 vssd1 vccd1 vccd1 _15390_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13354__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1779 _13984_/Q vssd1 vssd1 vccd1 vccd1 hold1779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _13671_/A1 hold2243/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07766_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ hold455/A hold549/A _14640_/Q _14736_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09506_/B sky130_fd_sc_hd__mux4_1
XANTENNA__08187__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09810__A2_N _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout634_A _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ hold537/X _13703_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold538/A sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09714_/A _09712_/B _09437_/C _09437_/D vssd1 vssd1 vccd1 vccd1 _09436_/X
+ sky130_fd_sc_hd__and4_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _14348_/Q _14252_/Q hold583/A _14124_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09368_/B sky130_fd_sc_hd__mux4_1
XANTENNA_fanout801_A _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07498__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08318_ _08318_/A _08318_/B _08318_/C vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__and3_1
XFILLER_0_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09298_ _08685_/C _10129_/A _09130_/X _09131_/X _10126_/A vssd1 vssd1 vccd1 vccd1
+ _09303_/A sky130_fd_sc_hd__a32o_1
XANTENNA_50 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 _11762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_72 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _07900_/B _08248_/Y _08208_/X vssd1 vssd1 vccd1 vccd1 _08250_/B sky130_fd_sc_hd__a21oi_4
XANTENNA_83 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_94 _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13545__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__C _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _11029_/X _11033_/C _11329_/B _11259_/X vssd1 vssd1 vccd1 vccd1 _11328_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_160_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10211_ _10386_/A _10209_/Y _09997_/B _10056_/A vssd1 vssd1 vccd1 vccd1 _10211_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11748__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _11620_/A _11614_/B vssd1 vssd1 vccd1 vccd1 _11192_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07775__A0 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ _10142_/A _10142_/B _14956_/Q _11623_/B vssd1 vssd1 vccd1 vccd1 _10312_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_207_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput190 _15171_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[6] sky130_fd_sc_hd__buf_12
XANTENNA__09516__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _10073_/A _10265_/A _10073_/C vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__and3_1
X_14950_ _15222_/CLK _14950_/D vssd1 vssd1 vccd1 vccd1 _14950_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12746__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ _15434_/CLK _13901_/D vssd1 vssd1 vccd1 vccd1 _13901_/Q sky130_fd_sc_hd__dfxtp_1
X_14881_ _14889_/CLK _14881_/D vssd1 vssd1 vccd1 vccd1 _14881_/Q sky130_fd_sc_hd__dfxtp_1
X_13832_ _15077_/CLK hold860/X vssd1 vssd1 vccd1 vccd1 hold859/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07262__A _15227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ hold179/X vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10975_ _10974_/B _10974_/C _10974_/A vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ hold2810/X _14218_/Q _14154_/Q hold1623/X _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12714_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_211_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13694_ hold199/X hold183/X _13698_/S vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15433_ _15433_/CLK _15433_/D vssd1 vssd1 vccd1 vccd1 _15433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12645_ _12645_/A _12645_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11512__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15364_ _15364_/CLK _15364_/D vssd1 vssd1 vccd1 vccd1 _15364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ _12601_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _12577_/C sky130_fd_sc_hd__or2_1
XFILLER_0_0_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07201__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ _15373_/CLK hold638/X vssd1 vssd1 vccd1 vccd1 hold637/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11527_ _11527_/A _11527_/B vssd1 vssd1 vccd1 vccd1 _11528_/B sky130_fd_sc_hd__xor2_1
X_15295_ _15424_/CLK _15295_/D vssd1 vssd1 vccd1 vccd1 _15295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14246_ _15372_/CLK _14246_/D vssd1 vssd1 vccd1 vccd1 _14246_/Q sky130_fd_sc_hd__dfxtp_1
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _11459_/A _11459_/B vssd1 vssd1 vccd1 vccd1 _11557_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11658__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13551__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _13584_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__nand2_1
X_14177_ _15179_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 _14177_/Q sky130_fd_sc_hd__dfxtp_1
X_11389_ _11588_/A _11623_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11390_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12343__A _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13491_/A hold137/X vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__and2_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13158__B _13158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ hold399/X _13924_/Q _13066_/S vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__mux2_1
Xhold1009 _14505_/Q vssd1 vssd1 vccd1 vccd1 hold1009/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12511__B1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09652__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13174__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ hold1391/X _13693_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13067__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07551_ _13386_/A hold175/X vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__and2_1
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08494__A1 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ hold1427/X _13721_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07482_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08494__B2 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _09494_/A1 _09094_/Y _09220_/X vssd1 vssd1 vccd1 vccd1 _09221_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13621__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12578__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _11333_/B _09709_/B _15210_/Q _08908_/A vssd1 vssd1 vccd1 vccd1 _09154_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08246__A1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09443__B1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__B2 _06939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08207__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12673__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07111__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ hold2758/X _08526_/B _12221_/B _08102_/Y _08100_/X vssd1 vssd1 vccd1 vccd1
+ _13379_/B sky130_fd_sc_hd__a221o_4
XFILLER_0_127_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11141__B _14970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13790__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09084_/B sky130_fd_sc_hd__or2_1
XFILLER_0_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08034_ _09918_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _08034_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput70 in0[14] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_1
XFILLER_0_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput81 in0[24] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_1
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12425__S0 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold810 hold810/A vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10980__B _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold821 hold821/A vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 in0[5] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_1
Xhold832 hold832/A vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_171_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold843 hold843/A vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13349__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 hold854/A vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 hold865/A vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 hold876/A vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 hold887/A vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 hold898/A vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _09984_/B _09984_/C _09984_/A vssd1 vssd1 vccd1 vccd1 _09987_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2200 _11760_/X vssd1 vssd1 vccd1 vccd1 _14554_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2211 _13920_/Q vssd1 vssd1 vccd1 vccd1 hold2211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08936_ _08933_/A _08934_/Y _08814_/B _08816_/B vssd1 vssd1 vccd1 vccd1 _08936_/Y
+ sky130_fd_sc_hd__o211ai_4
Xhold2222 _07455_/X vssd1 vssd1 vccd1 vccd1 _14085_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2233 _13953_/Q vssd1 vssd1 vccd1 vccd1 hold2233/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2244 _07766_/X vssd1 vssd1 vccd1 vccd1 _14382_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_186_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1510 _13520_/X vssd1 vssd1 vccd1 vccd1 _15278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2255 _13887_/Q vssd1 vssd1 vccd1 vccd1 hold2255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1521 _14758_/Q vssd1 vssd1 vccd1 vccd1 hold1521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2266 _11743_/X vssd1 vssd1 vccd1 vccd1 _14537_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2277 _13937_/Q vssd1 vssd1 vccd1 vccd1 hold2277/X sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ hold581/A _15275_/Q _15083_/Q _14376_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _08867_/X sky130_fd_sc_hd__mux4_1
Xhold1532 _07484_/X vssd1 vssd1 vccd1 vccd1 _14112_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2288 _07089_/X vssd1 vssd1 vccd1 vccd1 _13902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 _15435_/Q vssd1 vssd1 vccd1 vccd1 hold1543/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08182__B1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2299 _14912_/Q vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 _07730_/X vssd1 vssd1 vccd1 vccd1 _14349_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_66_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1565 _14475_/Q vssd1 vssd1 vccd1 vccd1 hold1565/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__B _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1576 _11966_/X vssd1 vssd1 vccd1 vccd1 _14785_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07818_ _12243_/A _07813_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _07818_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _08797_/A _08797_/B _08797_/C vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__a21oi_1
Xhold1587 _14303_/Q vssd1 vssd1 vccd1 vccd1 hold1587/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08178__A _08179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1598 _07605_/X vssd1 vssd1 vccd1 vccd1 _14229_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07749_ _13654_/A1 hold1209/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07749_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12805__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12900__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ _11493_/A _10757_/X _10759_/X vssd1 vssd1 vccd1 vccd1 _10760_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08906__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _09417_/B _09417_/C _09417_/A vssd1 vssd1 vccd1 vccd1 _09420_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10691_ _10691_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_165_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12430_ _12327_/A _12429_/X _12427_/X vssd1 vssd1 vccd1 vccd1 _13144_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13230__A1 _15062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12664__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12361_ _14268_/Q _14204_/Q _14140_/Q _14458_/Q _12365_/S0 _12343_/A vssd1 vssd1
+ vccd1 vccd1 _12361_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _14105_/CLK hold322/X vssd1 vssd1 vccd1 vccd1 _14100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11312_ _14296_/Q hold823/A hold357/A _14486_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _11313_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_133_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15080_ _15080_/CLK hold982/X vssd1 vssd1 vccd1 vccd1 hold981/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _15349_/Q _15348_/Q vssd1 vssd1 vccd1 vccd1 _13241_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_106_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_139_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14031_ _15199_/CLK _14031_/D vssd1 vssd1 vccd1 vccd1 _14031_/Q sky130_fd_sc_hd__dfxtp_1
X_11243_ _11620_/A _11564_/B _11000_/X _11001_/X _11542_/B vssd1 vssd1 vccd1 vccd1
+ _11248_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_28_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07257__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _11174_/A _11174_/B _11174_/C vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13693__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ _10296_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__and2_1
XANTENNA__13297__A1 input138/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07691__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10056_ _10056_/A _10056_/B _10056_/C _10056_/D vssd1 vssd1 vccd1 vccd1 _10056_/Y
+ sky130_fd_sc_hd__nand4_2
X_14933_ _15256_/CLK _14933_/D vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08173__B1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11507__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08088__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ _14866_/CLK _14864_/D vssd1 vssd1 vccd1 vccd1 _14864_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ _15276_/CLK _13815_/D vssd1 vssd1 vccd1 vccd1 _13815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14795_ _15441_/CLK hold640/X vssd1 vssd1 vccd1 vccd1 hold639/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11941__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13746_ hold829/X _13746_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold830/A sky130_fd_sc_hd__mux2_1
X_10958_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10958_/X sky130_fd_sc_hd__or2_1
XFILLER_0_128_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13441__B _13441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13677_ hold315/X hold2765/A _13682_/S vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__mux2_1
X_10889_ _10704_/B _10707_/B _10887_/X _10888_/Y vssd1 vssd1 vccd1 vccd1 _10889_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_183_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10784__C _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12628_ _13663_/A1 _12329_/B _12953_/B1 _13184_/B vssd1 vssd1 vccd1 vccd1 _12628_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15416_ _15416_/CLK hold820/X vssd1 vssd1 vccd1 vccd1 hold819/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09425__B1 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09976__A1 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15347_ _15424_/CLK _15347_/D vssd1 vssd1 vccd1 vccd1 _15347_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_182_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ hold765/X hold1729/X _12566_/S vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09647__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15278_ _15278_/CLK _15278_/D vssd1 vssd1 vccd1 vccd1 _15278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10008__D _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _14776_/CLK _14229_/D vssd1 vssd1 vccd1 vccd1 _14229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout608 _11407_/A vssd1 vssd1 vccd1 vccd1 _09858_/C sky130_fd_sc_hd__buf_8
XFILLER_0_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout619 _15205_/Q vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__10305__B _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _11473_/A _09764_/X _09766_/Y _09769_/X vssd1 vssd1 vccd1 vccd1 _13394_/B
+ sky130_fd_sc_hd__a31o_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13288__A1 input135/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06982_ _13654_/A1 hold1063/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06982_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12801__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08680_/X _08721_/B _08721_/C vssd1 vssd1 vccd1 vccd1 _08721_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_0_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ _15370_/Q _15273_/Q _15081_/Q _14374_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08652_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_178_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07603_ _11921_/A0 hold1457/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07603_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07106__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10678__D _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ _09661_/A _09712_/A vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__and2_1
XFILLER_0_194_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09113__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13632__A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07534_ hold389/X _13705_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold390/A sky130_fd_sc_hd__mux2_1
XFILLER_0_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08467__B2 _13182_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07465_ _13501_/A hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08562__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09204_ _09762_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__or2_1
XFILLER_0_147_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07396_ hold271/X _07450_/B vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__and2_1
XFILLER_0_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12646__S0 _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ _09136_/A _09253_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _09135_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__09511__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07776__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09066_ _09196_/A _09064_/C _08948_/B vssd1 vssd1 vccd1 vccd1 _09066_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08017_ _08091_/A _08017_/B _08017_/C vssd1 vssd1 vccd1 vccd1 _08091_/B sky130_fd_sc_hd__nand3_1
XANTENNA_fanout799_A _14490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12949__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 hold640/A vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13071__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold651 hold651/A vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 hold662/A vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold673 hold673/A vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 hold684/A vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 hold695/A vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13279__A1 input132/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__xnor2_2
Xhold2030 _07611_/X vssd1 vssd1 vccd1 vccd1 _14234_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2041 _14384_/Q vssd1 vssd1 vccd1 vccd1 hold2041/X sky130_fd_sc_hd__dlygate4sd3_1
X_08919_ _09164_/A _09676_/D _08920_/A vssd1 vssd1 vccd1 vccd1 _08919_/X sky130_fd_sc_hd__and3_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2052 _07762_/X vssd1 vssd1 vccd1 vccd1 _14378_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2063 _13903_/Q vssd1 vssd1 vccd1 vccd1 hold2063/X sky130_fd_sc_hd__dlygate4sd3_1
X_09899_ _09896_/Y _09897_/X _09742_/Y _09745_/X vssd1 vssd1 vccd1 vccd1 _09899_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2074 _13528_/X vssd1 vssd1 vccd1 vccd1 _15286_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1340 _07037_/X vssd1 vssd1 vccd1 vccd1 _13854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2085 _14235_/Q vssd1 vssd1 vccd1 vccd1 hold2085/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1351 _14786_/Q vssd1 vssd1 vccd1 vccd1 hold1351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2096 _07093_/X vssd1 vssd1 vccd1 vccd1 _13906_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11930_ _13718_/A1 hold1005/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11930_/X sky130_fd_sc_hd__mux2_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1362 _07162_/X vssd1 vssd1 vccd1 vccd1 _13970_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1373 _14379_/Q vssd1 vssd1 vccd1 vccd1 hold1373/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1384 _11813_/X vssd1 vssd1 vccd1 vccd1 _14637_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07016__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1395 _15441_/Q vssd1 vssd1 vccd1 vccd1 hold1395/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ hold469/X _13748_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold470/A sky130_fd_sc_hd__mux2_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13600_ input33/X _13634_/B _13625_/B vssd1 vssd1 vccd1 vccd1 _15326_/D sky130_fd_sc_hd__o21a_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11761__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10812_ _10812_/A _10978_/B _10812_/C vssd1 vssd1 vccd1 vccd1 _10814_/B sky130_fd_sc_hd__nand3_4
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13542__A _14427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _15408_/CLK hold270/X vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11057__A3 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ hold703/X _13679_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold704/A sky130_fd_sc_hd__mux2_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08636__A _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _13679_/A1 hold963/X _13534_/S vssd1 vssd1 vccd1 vccd1 hold964/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _10744_/A _10744_/B vssd1 vssd1 vccd1 vccd1 _10745_/A sky130_fd_sc_hd__or2_1
XANTENNA__11062__A _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13462_ _11106_/B _12288_/B _13468_/A vssd1 vssd1 vccd1 vccd1 _13463_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _10673_/A _10673_/B _10673_/C _10673_/D vssd1 vssd1 vccd1 vccd1 _10674_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _15324_/CLK _15201_/D vssd1 vssd1 vccd1 vccd1 _15201_/Q sky130_fd_sc_hd__dfxtp_4
X_12413_ _12642_/B1 _12408_/X _12412_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12420_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13688__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13754__A2 _12261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13393_ _13393_/A _13393_/B vssd1 vssd1 vccd1 vccd1 _15184_/D sky130_fd_sc_hd__and2_1
XFILLER_0_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11765__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15132_ _15132_/CLK _15132_/D vssd1 vssd1 vccd1 vccd1 _15132_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07686__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ hold1653/X hold1647/X _12466_/S vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15063_ _15063_/CLK _15063_/D vssd1 vssd1 vccd1 vccd1 _15063_/Q sky130_fd_sc_hd__dfxtp_1
X_12275_ _13487_/A _12275_/B vssd1 vssd1 vccd1 vccd1 _14924_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14014_ _15093_/CLK _14014_/D vssd1 vssd1 vccd1 vccd1 _14014_/Q sky130_fd_sc_hd__dfxtp_1
X_11226_ _11566_/A _15224_/Q _11224_/Y _11337_/A vssd1 vssd1 vccd1 vccd1 _11228_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11936__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _11156_/B _11435_/B _11156_/A vssd1 vssd1 vccd1 vccd1 _11158_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ _11578_/A _11577_/A _10108_/C _14963_/Q vssd1 vssd1 vccd1 vccd1 _10280_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11088_ _11089_/A _11089_/B _11089_/C vssd1 vssd1 vccd1 vccd1 _11273_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11237__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _10038_/B _10038_/C _10038_/A vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14916_ _15079_/CLK _14916_/D vssd1 vssd1 vccd1 vccd1 _14916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ _14975_/CLK _14847_/D vssd1 vssd1 vccd1 vccd1 _14847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11128__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13452__A _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08449__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778_ _15418_/CLK _14778_/D vssd1 vssd1 vccd1 vccd1 _14778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10256__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ hold955/X _13729_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 hold956/A sky130_fd_sc_hd__mux2_1
XANTENNA__12068__A _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ _09712_/A _09858_/A vssd1 vssd1 vccd1 vccd1 _08530_/A sky130_fd_sc_hd__and2_1
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07181_ _13748_/A1 hold1615/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07181_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07596__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09377__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12953__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2729_A _15170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10316__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11508__A1 _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12800__S0 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 _07182_/Y vssd1 vssd1 vccd1 vccd1 _07198_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__12181__A1 _12114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout416 _13716_/Y vssd1 vssd1 vccd1 vccd1 _13748_/S sky130_fd_sc_hd__buf_8
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11846__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout427 _11829_/Y vssd1 vssd1 vccd1 vccd1 _11845_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__08924__A2 _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout438 _07644_/Y vssd1 vssd1 vccd1 vccd1 _07676_/S sky130_fd_sc_hd__clkbuf_16
Xfanout449 _07981_/A vssd1 vssd1 vccd1 vccd1 _13570_/B sky130_fd_sc_hd__buf_4
X_09753_ _09749_/Y _09750_/X _09604_/Y _09606_/Y vssd1 vssd1 vccd1 vccd1 _09754_/C
+ sky130_fd_sc_hd__a211o_1
X_06965_ _14080_/Q _14079_/Q vssd1 vssd1 vccd1 vccd1 _06968_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12469__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08137__B1 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _08926_/A _09437_/A _08703_/C _08806_/A vssd1 vssd1 vccd1 vccd1 _08705_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09684_ _09684_/A _09684_/B _09684_/C vssd1 vssd1 vccd1 vccd1 _09684_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09262__D _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08635_ _08635_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _08636_/A sky130_fd_sc_hd__nor2_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11119__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13362__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10590__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08566_ _12252_/B _08566_/B vssd1 vssd1 vccd1 vccd1 _08566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08456__A _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07517_ hold751/X _13721_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 hold752/A sky130_fd_sc_hd__mux2_1
XFILLER_0_194_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08497_ _08496_/B _08600_/A _08496_/A vssd1 vssd1 vccd1 vccd1 _08498_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07448_ _07448_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14078_/D sky130_fd_sc_hd__and2_1
XFILLER_0_162_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08860__A1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07379_ _15341_/Q _07401_/A _14063_/Q _06908_/Y _07376_/X vssd1 vssd1 vccd1 vccd1
+ _07379_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09118_ _08841_/A _08838_/X _08840_/B vssd1 vssd1 vccd1 vccd1 _09119_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10390_ _10560_/A _10389_/C _10389_/A vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_115_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09049_ _09049_/A _09049_/B _09049_/C vssd1 vssd1 vccd1 vccd1 _09049_/X sky130_fd_sc_hd__and3_2
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09168__A2 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ hold2610/X hold2701/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09799__S0 _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 hold470/A vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 hold481/A vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08376__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _10826_/X _10829_/X _11008_/X _11010_/Y vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 hold492/A vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07254__B _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _13068_/A1 _12959_/X _12961_/X vssd1 vssd1 vccd1 vccd1 _12962_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 _07496_/X vssd1 vssd1 vccd1 vccd1 _14124_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__A1 _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _13668_/A1 hold1917/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__mux2_1
X_14701_ _15056_/CLK hold988/X vssd1 vssd1 vccd1 vccd1 hold987/A sky130_fd_sc_hd__dfxtp_1
Xhold1181 _14270_/Q vssd1 vssd1 vccd1 vccd1 hold1181/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__B2 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1192 _11774_/X vssd1 vssd1 vccd1 vccd1 _14599_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _13024_/S1 _12890_/X _12892_/X vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__a21o_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13272__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _15268_/CLK _14632_/D vssd1 vssd1 vccd1 vccd1 _14632_/Q sky130_fd_sc_hd__dfxtp_1
X_11844_ hold791/X hold2821/X _11845_/S vssd1 vssd1 vccd1 vccd1 hold792/A sky130_fd_sc_hd__mux2_1
XFILLER_0_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12858__S0 _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07270__A _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14563_ _14595_/CLK hold188/X vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ hold1189/X _13662_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10728_/B vssd1 vssd1 vccd1 vccd1 _10726_/Y sky130_fd_sc_hd__inv_2
X_13514_ _13662_/A1 hold705/X _13518_/S vssd1 vssd1 vccd1 vccd1 hold706/A sky130_fd_sc_hd__mux2_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14494_ _15428_/CLK _14494_/D vssd1 vssd1 vccd1 vccd1 _14494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13445_ _09625_/A _13450_/A _13444_/Y _13579_/C1 vssd1 vssd1 vccd1 vccd1 _15216_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ _11570_/A _11390_/A _10836_/A _10656_/D vssd1 vssd1 vccd1 vccd1 _10658_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13211__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10097__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ _13477_/A _13376_/B vssd1 vssd1 vccd1 vccd1 _15167_/D sky130_fd_sc_hd__and2_1
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10588_ _14292_/Q _14228_/Q _14164_/Q _14482_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _10589_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15115_ _15116_/CLK _15115_/D vssd1 vssd1 vccd1 vccd1 _15115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12327_ _12327_/A vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10961__A2 _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ _15270_/CLK _15046_/D vssd1 vssd1 vccd1 vccd1 _15046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _12254_/X _12257_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _13375_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12163__A1 hold2509/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11666__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _11209_/A _11209_/B _11209_/C vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12189_ hold2564/X _12195_/A2 _12188_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07445__A _08345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11674__A0 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08765__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08420_ _08420_/A _08516_/A _08420_/C vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__and3_1
XANTENNA__13182__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08276__A _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10229__A1 _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11414__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ _08352_/B _08441_/B _08350_/Y _13565_/C1 vssd1 vssd1 vccd1 vccd1 _08351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ _07302_/A _07302_/B vssd1 vssd1 vccd1 vccd1 _07319_/D sky130_fd_sc_hd__nand2_2
X_08282_ _08873_/A _08281_/X _08880_/A1 vssd1 vssd1 vccd1 vccd1 _08282_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07233_ _08169_/B _07233_/B vssd1 vssd1 vccd1 vccd1 _07323_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12526__A _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ _13665_/A1 hold1073/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07164_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07095_ _13698_/A1 hold2081/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07095_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12960__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout497_A _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13357__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__B1 _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _11320_/A _09805_/B vssd1 vssd1 vccd1 vccd1 _09805_/Y sky130_fd_sc_hd__nor2_1
X_07997_ _08065_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07997_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_157_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13103__B1 _12330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09736_ _09590_/Y _09592_/X _09734_/Y _09735_/X vssd1 vssd1 vccd1 vccd1 _09841_/A
+ sky130_fd_sc_hd__a211oi_1
X_06948_ _14027_/Q _14026_/Q _06953_/A vssd1 vssd1 vccd1 vccd1 _06950_/B sky130_fd_sc_hd__or3_1
Xclkbuf_4_12__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_88_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09667_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09667_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_179_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08756__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout831_A _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__A3 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _08617_/B _08617_/C _08617_/A vssd1 vssd1 vccd1 vccd1 _08618_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11605__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09598_ _09597_/B _09597_/C _09597_/A vssd1 vssd1 vccd1 vccd1 _09599_/C sky130_fd_sc_hd__a21oi_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08549_ _08201_/A _08548_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08549_/X sky130_fd_sc_hd__o21a_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _14947_/Q _11620_/B _11354_/B vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ _10510_/A _10510_/B _10510_/C vssd1 vssd1 vccd1 vccd1 _10513_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_162_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10640__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11491_ _13598_/A _11486_/Y _11490_/Y vssd1 vssd1 vccd1 vccd1 _11491_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12495__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11340__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12917__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ hold393/X _15062_/Q _13236_/S vssd1 vssd1 vccd1 vccd1 hold394/A sky130_fd_sc_hd__mux2_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _11577_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12393__A1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13161_ _13389_/A _13161_/B vssd1 vssd1 vccd1 vccd1 _15026_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10373_ _10373_/A _10373_/B _10373_/C vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__or3_2
X_12112_ _12112_/A _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12112_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ _13092_/A1 _13091_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12145__A1 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _12059_/A _12043_/B vssd1 vssd1 vccd1 vccd1 _14834_/D sky130_fd_sc_hd__and2_1
XANTENNA__07265__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10251__S0 _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 _11335_/A vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout791 _13076_/A vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__buf_6
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13645__A1 _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__B1 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ _15394_/CLK _13994_/D vssd1 vssd1 vccd1 vccd1 _13994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11656__A0 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12945_/A _12945_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _12952_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13206__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_140 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ _13101_/A _12876_/B vssd1 vssd1 vccd1 vccd1 _12877_/C sky130_fd_sc_hd__or2_1
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07204__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_151 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_162 _15007_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_173 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ _14791_/CLK _14615_/D vssd1 vssd1 vccd1 vccd1 _14615_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ hold341/X _13681_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold342/A sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _15411_/CLK _14546_/D vssd1 vssd1 vccd1 vccd1 _14546_/Q sky130_fd_sc_hd__dfxtp_1
X_11758_ _13711_/A1 hold869/X _11761_/S vssd1 vssd1 vccd1 vccd1 hold870/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _10532_/B _10534_/B _10706_/X _10708_/Y vssd1 vssd1 vccd1 vccd1 _10709_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11689_ input47/X _13648_/B vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__or2_1
X_14477_ _15411_/CLK _14477_/D vssd1 vssd1 vccd1 vccd1 _14477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13428_ _13440_/S _13428_/B vssd1 vssd1 vccd1 vccd1 _13428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13359_ _13360_/A _13359_/B vssd1 vssd1 vccd1 vccd1 _15150_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13008__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13333__B1 fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ _07920_/A _07920_/B vssd1 vssd1 vccd1 vccd1 _07921_/B sky130_fd_sc_hd__and2_1
X_15029_ _15190_/CLK _15029_/D vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dfxtp_1
Xhold2607 _14982_/Q vssd1 vssd1 vccd1 vccd1 hold2607/X sky130_fd_sc_hd__buf_2
Xhold2618 _12153_/X vssd1 vssd1 vccd1 vccd1 _14887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2629 _12141_/X vssd1 vssd1 vccd1 vccd1 _14881_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07851_ _07218_/X _07850_/X _07849_/X vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__a21oi_4
Xhold1906 _07596_/X vssd1 vssd1 vccd1 vccd1 _14220_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10242__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1917 _14734_/Q vssd1 vssd1 vccd1 vccd1 hold1917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1928 _11677_/X vssd1 vssd1 vccd1 vccd1 _14480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1939 _14788_/Q vssd1 vssd1 vccd1 vccd1 hold1939/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 dmemresp_rdata[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_07782_ hold381/X _13687_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold382/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ hold103/X _11514_/A2 _11514_/B1 _13191_/B _09519_/Y vssd1 vssd1 vccd1 vccd1
+ _09521_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09935__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12844__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__C _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11425__A _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12020__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ _09008_/A _08776_/A _08809_/D vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__and3_1
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11144__B _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09383_ _09816_/A _09809_/C vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08334_ _08240_/A _08240_/B _08242_/X vssd1 vssd1 vccd1 vccd1 _08335_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__13640__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10622__A1 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__C1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10622__B2 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ _08353_/B _08264_/Y _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08265_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout412_A _07080_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12256__A _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07216_ _07428_/A _07425_/A _07424_/A _07334_/C vssd1 vssd1 vccd1 vccd1 _09344_/B
+ sky130_fd_sc_hd__and4_4
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08196_ hold851/A _14241_/Q hold441/A _14113_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08197_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12375__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12690__S _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07147_ _13748_/A1 hold1343/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07147_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09240__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07784__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _14088_/Q _14089_/Q _14090_/Q vssd1 vssd1 vccd1 vccd1 _07115_/A sky130_fd_sc_hd__and3_2
XANTENNA_fanout781_A _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput350 _14817_/Q vssd1 vssd1 vccd1 vccd1 out2[4] sky130_fd_sc_hd__buf_12
XFILLER_0_140_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout879_A _06946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09284__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11350__A2 _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13088__C1 hold2774/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09719_ _09717_/X _09719_/B vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__and2b_1
X_10991_ _10990_/B _10990_/C _10990_/A vssd1 vssd1 vccd1 vccd1 _10992_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11102__A2 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ _13080_/A1 _12729_/X _12727_/X vssd1 vssd1 vccd1 vccd1 _13156_/B sky130_fd_sc_hd__a21oi_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07024__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__B _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12692_/A1 _12660_/X _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10861__B2 _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12865__S _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11612_ _11612_/A _11612_/B vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__xnor2_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13550__A _14431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14400_ _15428_/CLK _14400_/D vssd1 vssd1 vccd1 vccd1 _14400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12592_ _12642_/A1 _12591_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__a21o_1
X_15380_ _15380_/CLK hold552/X vssd1 vssd1 vccd1 vccd1 hold551/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11543_ _11390_/A _10356_/C _11420_/X _11449_/A vssd1 vssd1 vccd1 vccd1 _11545_/A
+ sky130_fd_sc_hd__a211oi_1
X_14331_ _15360_/CLK _14331_/D vssd1 vssd1 vccd1 vccd1 _14331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ _14485_/CLK hold668/X vssd1 vssd1 vccd1 vccd1 hold667/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11474_ hold2441/X _11474_/A2 _11324_/X _11325_/Y _11473_/X vssd1 vssd1 vccd1 vccd1
+ _11474_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_162_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13696__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ hold527/X _13659_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 hold528/A sky130_fd_sc_hd__mux2_1
X_10425_ _14291_/Q _14227_/Q hold477/A _14481_/Q _10425_/S0 _10425_/S1 vssd1 vssd1
+ vccd1 vccd1 _10426_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09231__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ _15190_/CLK hold156/X vssd1 vssd1 vccd1 vccd1 _14193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07694__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ _13381_/A _13144_/B vssd1 vssd1 vccd1 vccd1 _15009_/D sky130_fd_sc_hd__nor2_1
X_10356_ _11541_/A _11351_/B _10356_/C _11536_/B vssd1 vssd1 vccd1 vccd1 _10524_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09782__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _13071_/X _13072_/X _13074_/X _13073_/X _13100_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _13076_/B sky130_fd_sc_hd__mux4_1
X_10287_ _10287_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12213__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ hold2538/X hold2724/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output331_A _14829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11944__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13444__B _13444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A1 _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ _15372_/CLK _13977_/D vssd1 vssd1 vccd1 vccd1 _13977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12928_ _13708_/A1 _13103_/A2 _13078_/B1 _13196_/B vssd1 vssd1 vccd1 vccd1 _12928_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _15449_/Q _13916_/Q _13066_/S vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__mux2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12054__A0 _12120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13460__A _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14529_ _15394_/CLK _14529_/D vssd1 vssd1 vccd1 vccd1 _14529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ _08257_/C _08049_/Y _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08050_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10080__A2 _13396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07001_ _13739_/A1 hold1761/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07001_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12357__A1 _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2711_A _15184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ _08997_/B _08954_/B vssd1 vssd1 vccd1 vccd1 _08955_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12406__A1_N _07974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2404 _14861_/Q vssd1 vssd1 vccd1 vccd1 hold2404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2415 _15037_/Q vssd1 vssd1 vccd1 vccd1 hold2415/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07109__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__A2 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2426 _14864_/Q vssd1 vssd1 vccd1 vccd1 hold2426/X sky130_fd_sc_hd__dlygate4sd3_1
X_07903_ _07812_/A _09344_/B _07903_/C vssd1 vssd1 vccd1 vccd1 _07903_/Y sky130_fd_sc_hd__nand3b_2
Xhold2437 _14862_/Q vssd1 vssd1 vccd1 vccd1 hold2437/X sky130_fd_sc_hd__dlygate4sd3_1
X_08883_ hold2744/X input6/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13186_/B sky130_fd_sc_hd__mux2_2
Xhold1703 _14223_/Q vssd1 vssd1 vccd1 vccd1 hold1703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2448 _14852_/Q vssd1 vssd1 vccd1 vccd1 hold2448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2459 _14869_/Q vssd1 vssd1 vccd1 vccd1 hold2459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1714 _07752_/X vssd1 vssd1 vccd1 vccd1 _14368_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11332__A2 _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11854__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1725 _14910_/Q vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10766__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _12243_/A _07833_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _07834_/Y sky130_fd_sc_hd__o21ai_1
Xhold1736 _07785_/X vssd1 vssd1 vccd1 vccd1 _14400_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 _14125_/Q vssd1 vssd1 vccd1 vccd1 hold1747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 _13228_/X vssd1 vssd1 vccd1 vccd1 _15092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1769 _13845_/Q vssd1 vssd1 vccd1 vccd1 hold1769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07765_ _13736_/A1 hold1213/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11155__A _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09504_ hold695/A _15280_/Q _15088_/Q _14381_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09504_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ hold1071/X _13669_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 _07696_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09435_ _09435_/A _09571_/A _09714_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _09437_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12685__S _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_A _15203_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13370__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _10246_/A _09366_/B vssd1 vssd1 vccd1 vccd1 _09366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ _09164_/A _08685_/C _08317_/C _08317_/D vssd1 vssd1 vccd1 vccd1 _08318_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_145_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ _09297_/A _09297_/B vssd1 vssd1 vccd1 vccd1 _09305_/A sky130_fd_sc_hd__nand2_1
XANTENNA_40 _15013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_62 _13172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08248_ _13381_/B vssd1 vssd1 vccd1 vccd1 _08248_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_73 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_84 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_95 _15208_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08179_ _08179_/A _08179_/B vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11040__D _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10210_ _09997_/B _10056_/A _10386_/A _10209_/Y vssd1 vssd1 vccd1 vccd1 _10386_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _11564_/B _11189_/X _11188_/X vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10141_ _10141_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput180 _15191_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[26] sky130_fd_sc_hd__buf_12
XANTENNA__11308__C1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput191 _15172_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[7] sky130_fd_sc_hd__buf_12
XANTENNA__07019__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10072_ _09763_/A _09763_/B _10071_/X vssd1 vssd1 vccd1 vccd1 _10073_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11764__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ _15433_/CLK _13900_/D vssd1 vssd1 vccd1 vccd1 _13900_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10757__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ _14989_/CLK _14880_/D vssd1 vssd1 vccd1 vccd1 _14880_/Q sky130_fd_sc_hd__dfxtp_1
X_13831_ _15261_/CLK hold756/X vssd1 vssd1 vccd1 vccd1 hold755/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07262__B _14971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ _10974_/A _10974_/B _10974_/C vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__and3_1
X_13762_ hold187/X vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12713_ _12917_/B1 _12708_/X _12712_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12720_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13693_ hold711/X _13693_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 hold712/A sky130_fd_sc_hd__mux2_1
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12036__A0 _12102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15432_ _15432_/CLK hold662/X vssd1 vssd1 vccd1 vccd1 hold661/A sky130_fd_sc_hd__dfxtp_1
X_12644_ _12644_/A1 _12639_/X _12643_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12645_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08374__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12587__A1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15363_ _15432_/CLK hold894/X vssd1 vssd1 vccd1 vccd1 hold893/A sky130_fd_sc_hd__dfxtp_1
X_12575_ _12571_/X _12572_/X _12574_/X _12573_/X _12669_/A1 _12700_/S1 vssd1 vssd1
+ vccd1 vccd1 _12576_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10598__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14314_ _15190_/CLK _14314_/D vssd1 vssd1 vccd1 vccd1 _14314_/Q sky130_fd_sc_hd__dfxtp_1
X_11526_ _11526_/A _15225_/Q vssd1 vssd1 vccd1 vccd1 _11527_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15294_ _15424_/CLK _15294_/D vssd1 vssd1 vccd1 vccd1 _15294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11939__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _11457_/A _11457_/B vssd1 vssd1 vccd1 vccd1 _11459_/B sky130_fd_sc_hd__xnor2_1
X_14245_ _15438_/CLK hold974/X vssd1 vssd1 vccd1 vccd1 hold973/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10408_ _13750_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _10408_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ _15179_/CLK hold176/X vssd1 vssd1 vccd1 vccd1 _14176_/Q sky130_fd_sc_hd__dfxtp_1
X_11388_ _11623_/A _11537_/A _11623_/B _11588_/A vssd1 vssd1 vccd1 vccd1 _11390_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _10338_/B _10338_/C _10338_/D _11526_/A vssd1 vssd1 vccd1 vccd1 _10340_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13127_ _13489_/A hold39/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__and2_1
XANTENNA__10144__A _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ hold783/X hold1895/X hold655/X hold795/X _13066_/S _13068_/A1 vssd1 vssd1
+ vccd1 vccd1 _13058_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_175_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12511__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _12063_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _14817_/D sky130_fd_sc_hd__and2_1
XANTENNA__13455__A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__B _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13174__B _13174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07550_ _13386_/A hold215/X vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__and2_1
XFILLER_0_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07481_ hold1027/X _13687_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07481_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08494__A2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13190__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07599__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _09918_/A _12276_/B _13358_/B _08256_/A _09219_/Y vssd1 vssd1 vccd1 vccd1
+ _09220_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07900__B _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _09661_/A _09676_/D vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__and2_1
XANTENNA__12578__B2 _13182_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A1 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2759_A _15172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__B2 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ _08102_/A _08102_/B vssd1 vssd1 vccd1 vccd1 _08102_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12673__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11849__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _07900_/B _13378_/B hold2373/X vssd1 vssd1 vccd1 vccd1 _08033_/Y sky130_fd_sc_hd__a21oi_1
Xinput60 imemresp_data[5] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold800 hold800/A vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 in0[15] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold811 hold811/A vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 in0[25] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_1
XFILLER_0_130_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10980__C _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput93 in0[6] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__buf_1
XANTENNA__11002__A1 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold822 hold822/A vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold833 hold833/A vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 hold844/A vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold855 hold855/A vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 hold866/A vssd1 vssd1 vccd1 vccd1 hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold877 hold877/A vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold888 hold888/A vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _09984_/A _09984_/B _09984_/C vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__nand3_4
Xhold899 hold899/A vssd1 vssd1 vccd1 vccd1 hold899/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2201 _14733_/Q vssd1 vssd1 vccd1 vccd1 hold2201/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2212 _07107_/X vssd1 vssd1 vccd1 vccd1 _13920_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08935_ _08814_/B _08816_/B _08933_/A _08934_/Y vssd1 vssd1 vccd1 vccd1 _08935_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2223 _13963_/Q vssd1 vssd1 vccd1 vccd1 hold2223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2234 _07143_/X vssd1 vssd1 vccd1 vccd1 _13953_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout577_A _07448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 _07691_/X vssd1 vssd1 vccd1 vccd1 _14311_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2245 _13939_/Q vssd1 vssd1 vccd1 vccd1 hold2245/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1511 _15327_/Q vssd1 vssd1 vccd1 vccd1 _07423_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13365__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2256 _07071_/X vssd1 vssd1 vccd1 vccd1 _13887_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2267 _14768_/Q vssd1 vssd1 vccd1 vccd1 hold2267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _11938_/X vssd1 vssd1 vccd1 vccd1 _14758_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2278 _07127_/X vssd1 vssd1 vccd1 vccd1 _13937_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ _08981_/A _08863_/X _08865_/X vssd1 vssd1 vccd1 vccd1 _08866_/Y sky130_fd_sc_hd__o21ai_1
Xhold1533 _14711_/Q vssd1 vssd1 vccd1 vccd1 hold1533/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1544 _13725_/X vssd1 vssd1 vccd1 vccd1 _15435_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2289 hold2825/X vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__buf_1
Xhold1555 _14470_/Q vssd1 vssd1 vccd1 vccd1 hold1555/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1566 _11672_/X vssd1 vssd1 vccd1 vccd1 _14475_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07817_ _12233_/A _07817_/B vssd1 vssd1 vccd1 vccd1 _07817_/Y sky130_fd_sc_hd__nand2_1
X_08797_ _08797_/A _08797_/B _08797_/C vssd1 vssd1 vccd1 vccd1 _08799_/A sky130_fd_sc_hd__and3_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1577 _14802_/Q vssd1 vssd1 vccd1 vccd1 hold1577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1588 _07683_/X vssd1 vssd1 vccd1 vccd1 _14303_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1599 _14164_/Q vssd1 vssd1 vccd1 vccd1 hold1599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07748_ _13653_/A1 hold1359/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07748_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12361__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07679_ hold743/X _13652_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold744/A sky130_fd_sc_hd__mux2_1
XANTENNA__08906__B _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12018__A0 hold2607/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _09420_/B vssd1 vssd1 vccd1 vccd1 _09418_/Y sky130_fd_sc_hd__inv_2
X_10690_ _10691_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12569__A1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3__f_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ _09349_/A _09349_/B vssd1 vssd1 vccd1 vccd1 _13359_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08868__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12664__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ hold525/A hold327/A _14396_/Q hold517/A _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12360_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11759__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ _11507_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11311_/Y sky130_fd_sc_hd__nor2_1
X_12291_ _13171_/A _13468_/B vssd1 vssd1 vccd1 vccd1 _14940_/D sky130_fd_sc_hd__nor2_1
X_14030_ _14083_/CLK hold574/X vssd1 vssd1 vccd1 vccd1 _14030_/Q sky130_fd_sc_hd__dfxtp_1
X_11242_ _11242_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10427__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11173_ _11174_/A _11174_/B _11174_/C vssd1 vssd1 vccd1 vccd1 _11173_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _11580_/A _11594_/B _10328_/A _10123_/D vssd1 vssd1 vccd1 vccd1 _10125_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13275__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _10056_/A _10056_/B _10056_/C _10056_/D vssd1 vssd1 vccd1 vccd1 _10055_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_101_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14932_ _15258_/CLK _14932_/D vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__dfxtp_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08369__A _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08173__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__A _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2790 _15112_/Q vssd1 vssd1 vccd1 vccd1 _08631_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _14866_/CLK _14863_/D vssd1 vssd1 vccd1 vccd1 _14863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08088__B _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13814_ _14472_/CLK _13814_/D vssd1 vssd1 vccd1 vccd1 _13814_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12257__B1 hold2787/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14794_ _15371_/CLK hold786/X vssd1 vssd1 vccd1 vccd1 hold785/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13745_ hold575/X _13745_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold576/A sky130_fd_sc_hd__mux2_1
XFILLER_0_202_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10957_ _10956_/A _10956_/B _11640_/B1 vssd1 vssd1 vccd1 vccd1 _10957_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_196_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13214__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08881__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ hold1327/X _13742_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 _13676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10888_ _10887_/B _10887_/C _10887_/A vssd1 vssd1 vccd1 vccd1 _10888_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07212__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15415_ _15415_/CLK hold420/X vssd1 vssd1 vccd1 vccd1 hold419/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12627_ _13027_/A _12627_/B _12627_/C vssd1 vssd1 vccd1 vccd1 _12627_/X sky130_fd_sc_hd__and3_1
XFILLER_0_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09425__A1 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09425__B2 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09976__A2 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ _15348_/CLK _15346_/D vssd1 vssd1 vccd1 vccd1 _15346_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ hold199/X hold1983/X hold429/X hold2799/X _12566_/S _12368_/A vssd1 vssd1
+ vccd1 vccd1 _12558_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_170_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11669__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ _11509_/A _11509_/B vssd1 vssd1 vccd1 vccd1 _11509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15277_ _15374_/CLK _15277_/D vssd1 vssd1 vccd1 vccd1 _15277_/Q sky130_fd_sc_hd__dfxtp_1
X_12489_ _14273_/Q hold801/A _14145_/Q _14463_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12489_/X sky130_fd_sc_hd__mux4_1
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07448__A _07448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228_ _14775_/CLK _14228_/D vssd1 vssd1 vccd1 vccd1 _14228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14159_ _15411_/CLK hold390/X vssd1 vssd1 vccd1 vccd1 hold389/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout609 _15208_/Q vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _13653_/A1 hold2151/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06981_/X sky130_fd_sc_hd__mux2_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14__f_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13185__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _08716_/X _08718_/Y _08611_/Y _08613_/X vssd1 vssd1 vccd1 vccd1 _08721_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11299__A1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _08981_/A _08648_/X _08650_/X vssd1 vssd1 vccd1 vccd1 _08651_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_206_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07602_ _13741_/A1 hold2205/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07602_/X sky130_fd_sc_hd__mux2_1
X_08582_ _09816_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ hold515/X _13704_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold516/A sky130_fd_sc_hd__mux2_1
XFILLER_0_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13632__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08467__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ _12037_/A hold49/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__and2_1
XFILLER_0_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ _09762_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09203_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07395_ hold313/X _07450_/B vssd1 vssd1 vccd1 vccd1 hold314/A sky130_fd_sc_hd__and2_1
XFILLER_0_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12646__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _08776_/B _09714_/C _09864_/D _09136_/A vssd1 vssd1 vccd1 vccd1 _09138_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ _09065_/A vssd1 vssd1 vccd1 vccd1 _09199_/A sky130_fd_sc_hd__inv_2
XFILLER_0_115_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12264__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08016_ _10873_/A _15201_/Q vssd1 vssd1 vccd1 vccd1 _08017_/C sky130_fd_sc_hd__and2_1
XFILLER_0_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold630 hold630/A vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold641 hold641/A vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13071__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold652 hold652/A vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 hold663/A vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/A vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 hold685/A vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07792__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold696 hold696/A vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09573__A _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _14942_/Q _10338_/D vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout861_A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2020 _07131_/X vssd1 vssd1 vccd1 vccd1 _13941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2031 _13818_/Q vssd1 vssd1 vccd1 vccd1 hold2031/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2042 _07768_/X vssd1 vssd1 vccd1 vccd1 _14384_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08918_ _09164_/A _09676_/D vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__nand2_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2053 _15076_/Q vssd1 vssd1 vccd1 vccd1 hold2053/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12203__S _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ _09742_/Y _09745_/X _09896_/Y _09897_/X vssd1 vssd1 vccd1 vccd1 _09898_/Y
+ sky130_fd_sc_hd__a211oi_4
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _07090_/X vssd1 vssd1 vccd1 vccd1 _13903_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1330 _06993_/X vssd1 vssd1 vccd1 vccd1 _13812_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2075 _13936_/Q vssd1 vssd1 vccd1 vccd1 hold2075/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1341 _14594_/Q vssd1 vssd1 vccd1 vccd1 hold1341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2086 _07612_/X vssd1 vssd1 vccd1 vccd1 _14235_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1352 _11967_/X vssd1 vssd1 vccd1 vccd1 _14786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2097 _15081_/Q vssd1 vssd1 vccd1 vccd1 hold2097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _08849_/A _09344_/B vssd1 vssd1 vccd1 vccd1 _08851_/C sky130_fd_sc_hd__and2_1
XFILLER_0_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1363 _14771_/Q vssd1 vssd1 vccd1 vccd1 hold1363/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1374 _07763_/X vssd1 vssd1 vccd1 vccd1 _14379_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1385 _14696_/Q vssd1 vssd1 vccd1 vccd1 hold1385/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1396 _13731_/X vssd1 vssd1 vccd1 vccd1 _15441_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ hold487/X hold2817/X _11861_/S vssd1 vssd1 vccd1 vccd1 hold488/A sky130_fd_sc_hd__mux2_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10978_/A _10810_/C _10810_/A vssd1 vssd1 vccd1 vccd1 _10812_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13542__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ hold623/X _13711_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold624/A sky130_fd_sc_hd__mux2_1
XFILLER_0_196_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09655__A1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11057__A4 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13451__A2 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13034__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ _13711_/A1 hold1609/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10742_ _11288_/A1 _10741_/X _10598_/X vssd1 vssd1 vccd1 vccd1 _12286_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_211_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07032__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11062__B _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ _10673_/A _10673_/B _10673_/C _10673_/D vssd1 vssd1 vccd1 vccd1 _10673_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13461_ _10921_/B _13468_/A _13460_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 _13461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07967__S _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ _15324_/CLK _15200_/D vssd1 vssd1 vccd1 vccd1 _15200_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_180_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12412_ _12689_/S1 _12409_/X _12411_/X vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12411__B1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _13396_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _15183_/D sky130_fd_sc_hd__and2_1
XFILLER_0_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07969__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15131_ _15132_/CLK _15131_/D vssd1 vssd1 vccd1 vccd1 _15131_/Q sky130_fd_sc_hd__dfxtp_1
X_12343_ _12343_/A _12343_/B vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__and2_1
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15062_ _15062_/CLK _15062_/D vssd1 vssd1 vccd1 vccd1 _15062_/Q sky130_fd_sc_hd__dfxtp_1
X_12274_ _13150_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _14923_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ _11526_/A _11333_/B _15222_/Q _15223_/Q vssd1 vssd1 vccd1 vccd1 _11337_/A
+ sky130_fd_sc_hd__and4_1
X_14013_ _15408_/CLK hold840/X vssd1 vssd1 vccd1 vccd1 hold839/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12902__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11156_ _11156_/A _11156_/B _11435_/B vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13209__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ _13674_/A1 _11514_/A2 _11514_/B1 _13195_/B _10105_/Y vssd1 vssd1 vccd1 vccd1
+ _10107_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_207_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11087_ _11087_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _11089_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12478__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07207__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__B1 _09245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _10038_/A _10038_/B _10038_/C vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__nand3_1
X_14915_ _15391_/CLK _14915_/D vssd1 vssd1 vccd1 vccd1 _14915_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12573__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11237__B _15226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ _14992_/CLK _14846_/D vssd1 vssd1 vccd1 vccd1 _14846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11128__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13452__B _13452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14777_ _15418_/CLK _14777_/D vssd1 vssd1 vccd1 vccd1 _14777_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_170_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ hold563/X _13744_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 hold564/A sky130_fd_sc_hd__mux2_1
XFILLER_0_175_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ hold2033/X _13728_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_50_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13659_ hold2131/X _13659_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11205__A1 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_185_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07180_ _13681_/A1 hold1507/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07180_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12953__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ _15422_/CLK _15329_/D vssd1 vssd1 vccd1 vccd1 _15329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12953__B2 _13197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_65_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12705__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__A1 _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 _07182_/Y vssd1 vssd1 vccd1 vccd1 _07214_/S sky130_fd_sc_hd__clkbuf_16
X_09821_ _10351_/A _10338_/D vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__nand2_1
Xfanout417 _13698_/S vssd1 vssd1 vccd1 vccd1 _13714_/S sky130_fd_sc_hd__buf_8
Xfanout428 _11829_/Y vssd1 vssd1 vccd1 vccd1 _11861_/S sky130_fd_sc_hd__buf_8
Xfanout439 _07512_/Y vssd1 vssd1 vccd1 vccd1 _07528_/S sky130_fd_sc_hd__buf_12
XFILLER_0_193_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _09604_/Y _09606_/Y _09749_/Y _09750_/X vssd1 vssd1 vccd1 vccd1 _09754_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA_clkbuf_leaf_123_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06964_ _07744_/A _14089_/Q _14090_/Q vssd1 vssd1 vccd1 vccd1 _07182_/A sky130_fd_sc_hd__or3_4
XANTENNA__08137__A1 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__B2 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08703_ _08926_/A _09437_/A _08703_/C _08806_/A vssd1 vssd1 vccd1 vccd1 _08806_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12564__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _09684_/A _09684_/B _09684_/C vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07896__B1 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _07900_/B _13385_/B hold2733/X vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_90_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_138_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08550_/Y _08555_/Y _08564_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08566_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_178_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout442_A _07389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07516_ hold359/X _13687_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 hold360/A sky130_fd_sc_hd__mux2_1
X_08496_ _08496_/A _08496_/B _08600_/A vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07447_ _08535_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _14077_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_170_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08860__A2 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07378_ _15342_/Q _07402_/A _14061_/Q _07862_/A _07377_/X vssd1 vssd1 vccd1 vccd1
+ _07381_/C sky130_fd_sc_hd__o221a_1
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12944__A1 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09117_ _09117_/A _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09117_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10507__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09048_ _09047_/B _09047_/C _09047_/A vssd1 vssd1 vccd1 vccd1 _09049_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12157__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold460 hold460/A vssd1 vssd1 vccd1 vccd1 hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09799__S1 _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 hold471/A vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _11564_/A _11378_/C _11010_/C _11010_/D vssd1 vssd1 vccd1 vccd1 _11010_/Y
+ sky130_fd_sc_hd__nand4_1
Xhold482 hold482/A vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 hold493/A vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08376__B2 _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07027__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _13092_/A1 _12960_/X _13100_/S0 vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__a21o_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 _11945_/X vssd1 vssd1 vccd1 vccd1 _14765_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11772__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _15405_/CLK hold738/X vssd1 vssd1 vccd1 vccd1 hold737/A sky130_fd_sc_hd__dfxtp_1
Xhold1171 _15090_/Q vssd1 vssd1 vccd1 vccd1 hold1171/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _13519_/A0 hold2201/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11912_/X sky130_fd_sc_hd__mux2_1
Xhold1182 _07649_/X vssd1 vssd1 vccd1 vccd1 _14270_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10486__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _14673_/Q vssd1 vssd1 vccd1 vccd1 hold1193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ _13092_/A1 _12891_/X _14490_/Q vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__a21o_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _15079_/CLK _14631_/D vssd1 vssd1 vccd1 vccd1 _14631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ hold597/X _13730_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 hold598/A sky130_fd_sc_hd__mux2_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15190__D _15190_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12858__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07270__B _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _15042_/CLK hold264/X vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ hold1191/X _13661_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13699__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13513_ _13661_/A1 hold2149/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13513_/X sky130_fd_sc_hd__mux2_1
X_10725_ _10553_/B _10552_/Y _10723_/Y _10724_/X vssd1 vssd1 vccd1 vccd1 _10728_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_161_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _14731_/CLK sky130_fd_sc_hd__clkbuf_16
X_14493_ _15261_/CLK hold290/X vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07697__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13444_ _13450_/A _13444_/B vssd1 vssd1 vccd1 vccd1 _13444_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08382__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ _11570_/A _11390_/A _10836_/A _10656_/D vssd1 vssd1 vccd1 vccd1 _10836_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output194_A _06951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13375_ _13477_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _15166_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10097__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ _11507_/A _10587_/B vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15114_ _15116_/CLK _15114_/D vssd1 vssd1 vccd1 vccd1 _15114_/Q sky130_fd_sc_hd__dfxtp_1
X_12326_ _12326_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09239__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11947__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ _15045_/CLK _15045_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
X_12257_ _07894_/C _12256_/Y hold2787/X _08526_/B vssd1 vssd1 vccd1 vccd1 _12257_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12632__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _11207_/B _11386_/B _11207_/A vssd1 vssd1 vccd1 vccd1 _11209_/C sky130_fd_sc_hd__a21o_1
X_12188_ _14905_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__or2_1
XFILLER_0_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07445__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ hold2768/X input22/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13201_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12546__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09867__A1 _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11682__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08557__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14829_ _14866_/CLK _14829_/D vssd1 vssd1 vccd1 vccd1 _14829_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13182__B _13182_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13415__A2 _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12849__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08350_ _08265_/X _08349_/X _08441_/B vssd1 vssd1 vccd1 vccd1 _08350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11426__A1 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07301_ _15219_/Q _14963_/Q vssd1 vssd1 vccd1 vccd1 _07302_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08281_ _15398_/Q _14533_/Q hold815/A _14757_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08281_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_152_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15441_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07232_ _15201_/Q _11550_/A vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__A _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2741_A _15188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ _13664_/A1 hold1613/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07163_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07094_ _13730_/A1 hold2059/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07094_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11857__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13638__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08358__A1 _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10165__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A _07879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12261__B _12261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _09789_/Y _09794_/Y _09803_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09805_/B sky130_fd_sc_hd__a221o_1
XANTENNA__13639__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07996_ _14657_/Q _13930_/Q hold811/A _13898_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07997_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13103__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B2 _13203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _09734_/B _09734_/C _09734_/A vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__o21a_1
X_06947_ hold77/A hold127/A vssd1 vssd1 vccd1 vccd1 _06953_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_158_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13373__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09666_ _09666_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__A4 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ _08617_/A _08617_/B _08617_/C vssd1 vssd1 vccd1 vccd1 _08617_/Y sky130_fd_sc_hd__nor3_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11605__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09597_ _09597_/A _09597_/B _09597_/C vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout824_A _14488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08548_ _13873_/Q hold891/A hold687/A _13809_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08548_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08479_ _08908_/A _09026_/B _08702_/B _09437_/A vssd1 vssd1 vccd1 vccd1 _08480_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_163_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_143_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15457_/CLK sky130_fd_sc_hd__clkbuf_16
X_10510_ _10510_/A _10510_/B _10510_/C vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10640__A2 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11490_ _13598_/A _11486_/Y _10233_/A vssd1 vssd1 vccd1 vccd1 _11490_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12917__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ _14966_/Q _10273_/B _10440_/X vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11340__B _15226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10372_ _10373_/A _10373_/B _10373_/C vssd1 vssd1 vccd1 vccd1 _10372_/Y sky130_fd_sc_hd__nor3_1
X_13160_ _13389_/A _13160_/B vssd1 vssd1 vccd1 vccd1 _15025_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12111_ hold2465/X _12065_/Y _12110_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12111_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11767__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ _14361_/Q _14265_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13548__A _14430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08349__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ hold2605/X hold2700/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07546__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08349__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10251__S1 _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout770 _10700_/A vssd1 vssd1 vccd1 vccd1 _08926_/A sky130_fd_sc_hd__clkbuf_8
Xfanout781 _11335_/A vssd1 vssd1 vccd1 vccd1 _09661_/A sky130_fd_sc_hd__buf_4
Xfanout792 _13101_/A vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09849__A1 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13993_ _15361_/CLK hold682/X vssd1 vssd1 vccd1 vccd1 hold681/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09849__B2 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13645__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12944_ _12950_/S0 _12939_/X _12943_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12945_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10700__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12853__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07281__A _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _12871_/X _12872_/X _12874_/X _12873_/X _13100_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _12876_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_200_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14614_ _15382_/CLK hold486/X vssd1 vssd1 vccd1 vccd1 hold485/A sky130_fd_sc_hd__dfxtp_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _13444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ hold727/X _13680_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold728/A sky130_fd_sc_hd__mux2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_174 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_185 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_196 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12700__S0 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14545_ _15411_/CLK _14545_/D vssd1 vssd1 vccd1 vccd1 _14545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_134_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15452_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _13743_/A1 hold827/X _11761_/S vssd1 vssd1 vccd1 vccd1 hold828/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12627__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13222__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ _10707_/B _10707_/C _10707_/A vssd1 vssd1 vccd1 vccd1 _10708_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _15410_/CLK _14476_/D vssd1 vssd1 vccd1 vccd1 _14476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ _13241_/A _13792_/A2 _11687_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _14489_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13427_ _08535_/B _13440_/S _13426_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15207_/D
+ sky130_fd_sc_hd__o211a_1
X_10639_ _11620_/A _11378_/D _10639_/C _10639_/D vssd1 vssd1 vccd1 vccd1 _10641_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13360_/A _13358_/B vssd1 vssd1 vccd1 vccd1 _15149_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13008__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ _07375_/X _12379_/B _12330_/A vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ input71/X fanout1/X _13288_/X vssd1 vssd1 vccd1 vccd1 _13290_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13333__A1 input152/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15028_ _15190_/CLK _15028_/D vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13177__B _13177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2608 _12151_/X vssd1 vssd1 vccd1 vccd1 _14886_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2619 _14431_/Q vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07850_ hold313/A hold281/A hold255/A hold271/A vssd1 vssd1 vccd1 vccd1 _07850_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10242__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1907 _14136_/Q vssd1 vssd1 vccd1 vccd1 hold1907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1918 _11913_/X vssd1 vssd1 vccd1 vccd1 _14734_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1929 _14147_/Q vssd1 vssd1 vccd1 vccd1 hold1929/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07781_ hold1325/X _13719_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 _07781_/X sky130_fd_sc_hd__mux2_1
Xinput3 dmemresp_rdata[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_0_78_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09520_ hold2711/X input11/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13191_/B sky130_fd_sc_hd__mux2_2
XANTENNA__13193__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09935__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13095__C_N _13076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09451_/X sky130_fd_sc_hd__and2_1
XANTENNA__11425__B _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__D _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08402_ _08776_/B _08926_/A vssd1 vssd1 vccd1 vccd1 _08406_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09382_ _09291_/A _09290_/B _09290_/A vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _08335_/B vssd1 vssd1 vccd1 vccd1 _08333_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_125_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15056_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08264_ _08352_/B _08352_/C vssd1 vssd1 vccd1 vccd1 _08264_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10622__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07130__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07215_ _15330_/Q _15327_/Q _15326_/Q _15331_/Q vssd1 vssd1 vccd1 vccd1 _07334_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08195_ _08760_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout405_A _07182_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09846__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _13714_/A1 hold1479/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07146_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13368__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__B _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ _13748_/A1 hold1817/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07077_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12272__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput340 _14837_/Q vssd1 vssd1 vccd1 vccd1 out2[24] sky130_fd_sc_hd__buf_12
XANTENNA__13324__A1 input148/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput351 _14818_/Q vssd1 vssd1 vccd1 vccd1 out2[5] sky130_fd_sc_hd__buf_12
XANTENNA__12127__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12758__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09284__C _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout774_A _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09581__A _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _08042_/B _14426_/Q vssd1 vssd1 vccd1 vccd1 _07979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09718_ _09715_/Y _09716_/X _09570_/X _09572_/X vssd1 vssd1 vccd1 vccd1 _09719_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10520__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10992_/B sky130_fd_sc_hd__nand3_2
XANTENNA__08197__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07937__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11335__B _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09649_ _10244_/A _09648_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09649_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_195_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__A2 _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ hold791/A _13940_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_210_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08925__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09520__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__xnor2_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12591_ hold631/A hold973/A _12591_/S vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_116_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15376_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11351__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14330_ _15390_/CLK _14330_/D vssd1 vssd1 vccd1 vccd1 _14330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11542_ _11542_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _11546_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07040__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _15454_/CLK hold904/X vssd1 vssd1 vccd1 vccd1 hold903/A sky130_fd_sc_hd__dfxtp_1
X_11473_ _11473_/A _11473_/B _11473_/C vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__and3_1
XFILLER_0_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ hold2053/X _13724_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10424_ _11493_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10424_/Y sky130_fd_sc_hd__nor2_1
X_14192_ _15188_/CLK hold194/X vssd1 vssd1 vccd1 vccd1 _14192_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08660__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13278__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ _13381_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _15008_/D sky130_fd_sc_hd__nor2_1
X_10355_ _10129_/A _10827_/D _10127_/X _10126_/X _11588_/A vssd1 vssd1 vccd1 vccd1
+ _10360_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13315__A1 input145/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07276__A _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12749__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ _11573_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__and2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _13892_/Q hold401/A _13860_/Q _13828_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux4_1
X_12025_ _12059_/A _12025_/B vssd1 vssd1 vccd1 vccd1 _14825_/D sky130_fd_sc_hd__and2_1
XFILLER_0_139_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08742__A1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13618__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13217__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11526__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ _15374_/CLK _13976_/D vssd1 vssd1 vccd1 vccd1 _13976_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09298__A2 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12921__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ _13102_/A _12927_/B _12927_/C vssd1 vssd1 vccd1 vccd1 _12927_/X sky130_fd_sc_hd__and3_1
XFILLER_0_198_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__S _11960_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ _15412_/Q _14547_/Q hold491/A _14771_/Q _13066_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12858_/X sky130_fd_sc_hd__mux4_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11809_ hold1227/X _13663_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11809_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13460__B _13460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_107_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _14889_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12789_ _14285_/Q _14221_/Q hold417/A _14475_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12789_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _15397_/CLK _14528_/D vssd1 vssd1 vccd1 vccd1 _14528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14459_ _15361_/CLK _14459_/D vssd1 vssd1 vccd1 vccd1 _14459_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12791__S _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07000_ _13705_/A1 hold1495/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13188__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12092__A _14986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13306__A1 input142/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ _08997_/A _08950_/C _08950_/A vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11317__B1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2405 _12099_/X vssd1 vssd1 vccd1 vccd1 _14861_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ _13653_/A1 _12260_/A2 _07901_/X _07882_/Y vssd1 vssd1 vccd1 vccd1 _12262_/B
+ sky130_fd_sc_hd__a211o_2
Xhold2416 _13749_/B vssd1 vssd1 vccd1 vccd1 _13406_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2427 _12105_/X vssd1 vssd1 vccd1 vccd1 _14864_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08882_ _11320_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08882_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_209_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2438 _12101_/X vssd1 vssd1 vccd1 vccd1 _14862_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08194__C1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1704 _07599_/X vssd1 vssd1 vccd1 vccd1 _14223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2449 _12081_/X vssd1 vssd1 vccd1 vccd1 _14852_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1715 _14772_/Q vssd1 vssd1 vccd1 vccd1 hold1715/X sky130_fd_sc_hd__dlygate4sd3_1
X_07833_ _15392_/Q _14527_/Q _14687_/Q _14751_/Q _12198_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _07833_/X sky130_fd_sc_hd__mux4_1
Xhold1726 _13471_/X vssd1 vssd1 vccd1 vccd1 _15230_/D sky130_fd_sc_hd__buf_1
Xhold1737 _14737_/Q vssd1 vssd1 vccd1 vccd1 hold1737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1748 _07497_/X vssd1 vssd1 vccd1 vccd1 _14125_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1759 _13798_/Q vssd1 vssd1 vccd1 vccd1 hold1759/X sky130_fd_sc_hd__dlygate4sd3_1
X_07764_ _13669_/A1 hold2119/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07764_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12817__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07125__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _09941_/A _09500_/X _09502_/X vssd1 vssd1 vccd1 vccd1 _09503_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11155__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12966__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07695_ hold637/X _13668_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold638/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11870__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09434_ _09435_/A _09571_/A _09714_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09434_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09365_ _10426_/A _09362_/X _09364_/X _10255_/A1 vssd1 vssd1 vccd1 vccd1 _09366_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout522_A _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ _09164_/A _08685_/C _08317_/C _08317_/D vssd1 vssd1 vccd1 vccd1 _08318_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ _09143_/A _09142_/B _09140_/X vssd1 vssd1 vccd1 vccd1 _09307_/A sky130_fd_sc_hd__a21o_1
XANTENNA_30 _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_41 _15013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 _12294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08247_ _12258_/S _08244_/X _08245_/Y _08246_/X vssd1 vssd1 vccd1 vccd1 _13381_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_74 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_85 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10359__A1 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08178_ _08179_/A _08179_/B vssd1 vssd1 vccd1 vccd1 _08178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout891_A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07129_ _13730_/A1 hold2245/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07129_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08972__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput170 _15182_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[17] sky130_fd_sc_hd__buf_12
XFILLER_0_98_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput181 _15192_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[27] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput192 _15173_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[8] sky130_fd_sc_hd__buf_12
X_10071_ _10071_/A _10071_/B _09766_/A vssd1 vssd1 vccd1 vccd1 _10071_/X sky130_fd_sc_hd__or3b_1
XANTENNA__11859__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _15296_/CLK _13830_/D vssd1 vssd1 vccd1 vccd1 _13830_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10250__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07035__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13761_ hold263/X vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _10972_/B _10972_/C _10972_/A vssd1 vssd1 vccd1 vccd1 _10974_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11780__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ _12749_/S1 _12709_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_167_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ hold1323/X hold285/X _13698_/S vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_195_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ _15433_/CLK hold812/X vssd1 vssd1 vccd1 vccd1 hold811/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12643_ _12699_/S1 _12640_/X _12642_/X vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_26_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ _15397_/CLK hold950/X vssd1 vssd1 vccd1 vccd1 hold949/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _13872_/Q _14000_/Q _13840_/Q _13808_/Q _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12574_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_142_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10598__B2 _13198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14313_ _15179_/CLK _14313_/D vssd1 vssd1 vccd1 vccd1 _14313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11525_ _11461_/A _11461_/B _11462_/Y vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__o21a_1
X_15293_ _15293_/CLK _15293_/D vssd1 vssd1 vccd1 vccd1 _15293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14244_ _14956_/CLK hold832/X vssd1 vssd1 vccd1 vccd1 hold831/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ _11457_/B _11457_/A vssd1 vssd1 vccd1 vccd1 _11557_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12744__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10407_ _11108_/A _10746_/A vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14175_ _15177_/CLK hold216/X vssd1 vssd1 vccd1 vccd1 _14175_/Q sky130_fd_sc_hd__dfxtp_1
X_11387_ _11168_/A _11588_/B _11165_/X _11166_/X _11606_/B vssd1 vssd1 vccd1 vccd1
+ _11392_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_22_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08963__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ _13129_/A hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__and2_1
X_10338_ _11526_/A _10338_/B _10338_/C _10338_/D vssd1 vssd1 vccd1 vccd1 _10338_/X
+ sky130_fd_sc_hd__and4_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11955__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13107_/A _13057_/B vssd1 vssd1 vccd1 vccd1 _14970_/D sky130_fd_sc_hd__nor2_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _10177_/A _10177_/B _10179_/X vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__a21oi_1
X_12008_ hold2628/X hold2671/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10798__C _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__B _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13959_ _15299_/CLK _13959_/D vssd1 vssd1 vccd1 vccd1 _13959_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13471__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07480_ hold517/X _13719_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 hold518/A sky130_fd_sc_hd__mux2_1
XFILLER_0_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07151__A0 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09150_ _09816_/A _09979_/C vssd1 vssd1 vccd1 vccd1 _09160_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12578__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09443__A2 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _07323_/C _08029_/X _08169_/B vssd1 vssd1 vccd1 vccd1 _08102_/B sky130_fd_sc_hd__a21oi_1
X_09081_ hold2569/X _09344_/B _09346_/B vssd1 vssd1 vccd1 vccd1 _09083_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13410__S _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09396__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ hold2648/X _08526_/B _08028_/X _08031_/X vssd1 vssd1 vccd1 vccd1 _13378_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_0_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 imemresp_data[25] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_1
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput61 imemresp_data[6] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput72 in0[16] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold801 hold801/A vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 hold812/A vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 in0[26] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold823 hold823/A vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 in0[7] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_1
XFILLER_0_130_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 hold834/A vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12026__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold845 hold845/A vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 hold856/A vssd1 vssd1 vccd1 vccd1 hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold878 hold878/A vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _09982_/B _10182_/B _09982_/A vssd1 vssd1 vccd1 vccd1 _09984_/C sky130_fd_sc_hd__a21o_1
Xhold889 hold889/A vssd1 vssd1 vccd1 vccd1 hold889/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11865__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2202 _11912_/X vssd1 vssd1 vccd1 vccd1 _14733_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ _08932_/B _08932_/C _08932_/A vssd1 vssd1 vccd1 vccd1 _08934_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__13646__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2213 _14420_/Q vssd1 vssd1 vccd1 vccd1 hold2213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2224 _07155_/X vssd1 vssd1 vccd1 vccd1 _13963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2235 _13825_/Q vssd1 vssd1 vccd1 vccd1 hold2235/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1501 _14538_/Q vssd1 vssd1 vccd1 vccd1 hold1501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2246 _07129_/X vssd1 vssd1 vccd1 vccd1 _13939_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1512 _07423_/X vssd1 vssd1 vccd1 vccd1 _14053_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08865_ _08989_/A _08864_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08865_/X sky130_fd_sc_hd__o21a_1
Xhold2257 _13958_/Q vssd1 vssd1 vccd1 vccd1 hold2257/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout472_A _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2268 _11948_/X vssd1 vssd1 vccd1 vccd1 _14768_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1523 _13968_/Q vssd1 vssd1 vccd1 vccd1 hold1523/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2279 _13919_/Q vssd1 vssd1 vccd1 vccd1 hold2279/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _11889_/X vssd1 vssd1 vccd1 vccd1 _14711_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11166__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1545 _14596_/Q vssd1 vssd1 vccd1 vccd1 hold1545/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08182__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1556 _11667_/X vssd1 vssd1 vccd1 vccd1 _14470_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07816_ _13864_/Q _13992_/Q _07816_/S vssd1 vssd1 vccd1 vccd1 _07817_/B sky130_fd_sc_hd__mux2_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1567 _14464_/Q vssd1 vssd1 vccd1 vccd1 hold1567/X sky130_fd_sc_hd__dlygate4sd3_1
X_08796_ _08686_/A _08686_/B _08686_/C vssd1 vssd1 vccd1 vccd1 _08797_/C sky130_fd_sc_hd__a21bo_1
Xhold1578 _11983_/X vssd1 vssd1 vccd1 vccd1 _14802_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 _14603_/Q vssd1 vssd1 vccd1 vccd1 hold1589/X sky130_fd_sc_hd__dlygate4sd3_1
X_07747_ _13652_/A1 hold2141/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07747_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout737_A _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13381__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12361__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ hold529/X _13651_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold530/A sky130_fd_sc_hd__mux2_1
XFILLER_0_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09417_ _09417_/A _09417_/B _09417_/C vssd1 vssd1 vccd1 vccd1 _09420_/B sky130_fd_sc_hd__and3_1
XFILLER_0_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ _09217_/A _09217_/B _09215_/A vssd1 vssd1 vccd1 vccd1 _09349_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08868__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09279_ _09459_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ hold657/A _14264_/Q hold473/A _14136_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _11311_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ _13107_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _14939_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11241_ _11014_/A _11013_/B _11011_/X vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10427__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11172_ _11563_/A _11605_/B vssd1 vssd1 vccd1 vccd1 _11174_/C sky130_fd_sc_hd__and2_1
XANTENNA__11775__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _11580_/A _14964_/Q _10328_/A _10123_/D vssd1 vssd1 vccd1 vccd1 _10296_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13556__A _14434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10054_ _10164_/A _10052_/C _10052_/A vssd1 vssd1 vccd1 vccd1 _10056_/D sky130_fd_sc_hd__a21o_1
XANTENNA__07554__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ _15244_/CLK _14931_/D vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2780 _11287_/X vssd1 vssd1 vccd1 vccd1 _13403_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2791 _15122_/Q vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07273__B _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ _14866_/CLK _14862_/D vssd1 vssd1 vccd1 vccd1 _14862_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13813_ _14409_/CLK _13813_/D vssd1 vssd1 vccd1 vccd1 _13813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13454__A0 _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__B2 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14793_ _15440_/CLK _14793_/D vssd1 vssd1 vccd1 vccd1 _14793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09122__A1 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ hold715/X _13744_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold716/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ hold843/X _13675_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold844/A sky130_fd_sc_hd__mux2_1
X_10887_ _10887_/A _10887_/B _10887_/C vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__and3_2
XFILLER_0_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _15451_/CLK _15414_/D vssd1 vssd1 vccd1 vccd1 _15414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _12676_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12627_/C sky130_fd_sc_hd__or2_1
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09425__A2 _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15345_ _15422_/CLK _15345_/D vssd1 vssd1 vccd1 vccd1 _15345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12607_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _14950_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09976__A3 _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13230__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10440__B1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _11504_/A _11505_/X _11507_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _11509_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_112_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15276_ _15276_/CLK hold948/X vssd1 vssd1 vccd1 vccd1 hold947/A sky130_fd_sc_hd__dfxtp_1
X_12488_ _12642_/B1 _12483_/X _12487_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12495_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ _15415_/CLK _14227_/D vssd1 vssd1 vccd1 vccd1 _14227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11439_ _11573_/A _11594_/B _11439_/C _11439_/D vssd1 vssd1 vccd1 vccd1 _11441_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__10418__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ _15410_/CLK hold516/X vssd1 vssd1 vccd1 vccd1 hold515/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13466__A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ _13495_/A hold159/X vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__and2_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14089_ _15214_/CLK _14089_/D vssd1 vssd1 vccd1 vccd1 _14089_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _13652_/A1 hold2217/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06980_/X sky130_fd_sc_hd__mux2_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09361__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08650_ _08989_/A _08649_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08650_/X sky130_fd_sc_hd__o21a_1
X_07601_ _13740_/A1 hold1293/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07601_/X sky130_fd_sc_hd__mux2_1
X_08581_ _08581_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07532_ hold417/X _13703_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold418/A sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07463_ hold273/X _13535_/B vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__and2_1
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09202_ _09202_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ hold281/X _07450_/B vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__and2_1
XFILLER_0_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09133_ _09133_/A _09133_/B vssd1 vssd1 vccd1 vccd1 _09143_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_115_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09064_ _08948_/B _09196_/A _09064_/C vssd1 vssd1 vccd1 vccd1 _09065_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08015_ _08014_/B _08014_/C _08014_/A vssd1 vssd1 vccd1 vccd1 _08017_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_170_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold620 hold620/A vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold631 hold631/A vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08927__A1 _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 hold642/A vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 hold653/A vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold664 hold664/A vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold675 hold675/A vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 hold686/A vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold697 hold697/A vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13376__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14910__D _14910_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12280__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2010 _11924_/X vssd1 vssd1 vccd1 vccd1 _14745_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2021 _13843_/Q vssd1 vssd1 vccd1 vccd1 hold2021/X sky130_fd_sc_hd__dlygate4sd3_1
X_08917_ _08917_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__xnor2_2
Xhold2032 _06999_/X vssd1 vssd1 vccd1 vccd1 _13818_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12487__A1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2043 _14129_/Q vssd1 vssd1 vccd1 vccd1 hold2043/X sky130_fd_sc_hd__dlygate4sd3_1
X_09897_ _09896_/A _09896_/B _09896_/C _09896_/D vssd1 vssd1 vccd1 vccd1 _09897_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2054 _13212_/X vssd1 vssd1 vccd1 vccd1 _15076_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _07165_/X vssd1 vssd1 vccd1 vccd1 _13973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2065 _14643_/Q vssd1 vssd1 vccd1 vccd1 hold2065/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15248_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _15387_/Q vssd1 vssd1 vccd1 vccd1 hold1331/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2076 _07126_/X vssd1 vssd1 vccd1 vccd1 _13936_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2087 _14729_/Q vssd1 vssd1 vccd1 vccd1 hold2087/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 _11769_/X vssd1 vssd1 vccd1 vccd1 _14594_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08848_ _07900_/B _13387_/B _08773_/X vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__a21o_4
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1353 _14722_/Q vssd1 vssd1 vccd1 vccd1 hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2098 _13217_/X vssd1 vssd1 vccd1 vccd1 _15081_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1364 _11951_/X vssd1 vssd1 vccd1 vccd1 _14771_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1375 _14503_/Q vssd1 vssd1 vccd1 vccd1 hold1375/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07902__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1386 _11874_/X vssd1 vssd1 vccd1 vccd1 _14696_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12239__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _08892_/A _09864_/C _09864_/D _08901_/A vssd1 vssd1 vccd1 vccd1 _08783_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 _14606_/Q vssd1 vssd1 vccd1 vccd1 hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ _10810_/A _10978_/A _10810_/C vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__nand3_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ hold1245/X hold2765/A _11795_/S vssd1 vssd1 vccd1 vccd1 _11790_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09655__A2 _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ hold2706/X _11474_/A2 _10602_/X _10740_/Y _10739_/Y vssd1 vssd1 vccd1 vccd1
+ _10741_/X sky130_fd_sc_hd__a221o_2
XANTENNA__07666__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13460_ _13468_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10672_ _10669_/A _10670_/Y _10496_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10673_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _12642_/A1 _12410_/X _12644_/A1 vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_152_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13391_ _13393_/A _13391_/B vssd1 vssd1 vccd1 vccd1 _15182_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12411__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15390_/CLK sky130_fd_sc_hd__clkbuf_16
X_15130_ _15132_/CLK _15130_/D vssd1 vssd1 vccd1 vccd1 _15130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07969__A2 _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ hold755/A _13799_/Q _12466_/S vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15061_ _15377_/CLK _15061_/D vssd1 vssd1 vccd1 vccd1 _15061_/Q sky130_fd_sc_hd__dfxtp_1
X_12273_ _13487_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _14922_/D sky130_fd_sc_hd__and2_1
XFILLER_0_65_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14012_ _15191_/CLK hold676/X vssd1 vssd1 vccd1 vccd1 hold675/A sky130_fd_sc_hd__dfxtp_1
X_11224_ _11333_/B _15222_/Q _15223_/Q _11526_/A vssd1 vssd1 vccd1 vccd1 _11224_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ _11590_/A _11594_/B _11155_/C _11435_/A vssd1 vssd1 vccd1 vccd1 _11435_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_207_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07284__A _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ hold2741/X input16/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13195_/B sky130_fd_sc_hd__mux2_2
X_11086_ _11086_/A _11086_/B _11087_/B vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__and3_1
XANTENNA__12478__B2 _13178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15387_/CLK sky130_fd_sc_hd__clkbuf_16
X_10037_ _10036_/B _10141_/B _10036_/A vssd1 vssd1 vccd1 vccd1 _10038_/C sky130_fd_sc_hd__a21o_1
X_14914_ _15367_/CLK _14914_/D vssd1 vssd1 vccd1 vccd1 _14914_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12573__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14845_ _14975_/CLK _14845_/D vssd1 vssd1 vccd1 vccd1 _14845_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13225__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07106__A0 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14776_ _14776_/CLK hold774/X vssd1 vssd1 vccd1 vccd1 hold773/A sky130_fd_sc_hd__dfxtp_1
X_11988_ hold1185/X hold2765/A _11993_/S vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13727_ hold765/X _13727_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 hold766/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10939_ _11493_/A _10939_/B vssd1 vssd1 vccd1 vccd1 _10939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ hold647/X _13724_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold648/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12938__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ hold955/A _13906_/Q _12641_/S vssd1 vssd1 vccd1 vccd1 _12609_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11205__A2 _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13589_ _10744_/B _13591_/A2 _13588_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _15320_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15316_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15328_ _15422_/CLK _15328_/D vssd1 vssd1 vccd1 vccd1 _15328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12953__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ _15389_/CLK hold114/X vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08385__A2 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _07149_/X vssd1 vssd1 vccd1 vccd1 _07165_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold2617_A _14983_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout418 _13715_/S vssd1 vssd1 vccd1 vccd1 _13698_/S sky130_fd_sc_hd__buf_12
XFILLER_0_120_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07593__A0 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 _11796_/Y vssd1 vssd1 vccd1 vccd1 _11812_/S sky130_fd_sc_hd__buf_12
X_09751_ _09604_/Y _09606_/Y _09749_/Y _09750_/X vssd1 vssd1 vccd1 vccd1 _09751_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11428__B _14971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06963_ _14027_/Q _06953_/A _06962_/X _06959_/X vssd1 vssd1 vccd1 vccd1 _06963_/X
+ sky130_fd_sc_hd__o31a_4
XANTENNA__12469__A1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15421_/CLK sky130_fd_sc_hd__clkbuf_16
X_08702_ _09138_/A _08702_/B _08809_/B _08809_/D vssd1 vssd1 vccd1 vccd1 _08806_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08137__A2 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09682_ _09681_/B _09681_/C _09681_/A vssd1 vssd1 vccd1 vccd1 _09684_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12564__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08633_ _12221_/B _08569_/X _08570_/Y _08632_/X vssd1 vssd1 vccd1 vccd1 _13385_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__07922__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11692__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08564_/A1 _08557_/Y _08559_/Y _08561_/Y _08563_/Y vssd1 vssd1 vccd1 vccd1
+ _08564_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07133__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07515_ hold2105/X _13719_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07515_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07648__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08495_ _08776_/A _08776_/B _08809_/B _08809_/D vssd1 vssd1 vccd1 vccd1 _08600_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout435_A _07710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ _08435_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _14076_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07377_ _07862_/C _14059_/Q _07403_/A _15343_/Q vssd1 vssd1 vccd1 vccd1 _07377_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout602_A _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12275__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ _13519_/A0 _11514_/A2 _11514_/B1 _13188_/B _09114_/Y vssd1 vssd1 vccd1 vccd1
+ _09116_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10507__B _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09047_ _09047_/A _09047_/B _09047_/C vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_62_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold450 hold450/A vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold461/A vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 hold472/A vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08376__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold483 hold483/A vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 hold494/A vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _11497_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _09949_/Y sky130_fd_sc_hd__nor2_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _14485_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ hold1673/X hold1571/X _13066_/S vssd1 vssd1 vccd1 vccd1 _12960_/X sky130_fd_sc_hd__mux2_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 _11755_/X vssd1 vssd1 vccd1 vccd1 _14549_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07832__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _13666_/A1 hold1407/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11911_/X sky130_fd_sc_hd__mux2_1
Xhold1161 _14275_/Q vssd1 vssd1 vccd1 vccd1 hold1161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 _13226_/X vssd1 vssd1 vccd1 vccd1 _15090_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12880__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ _14353_/Q _14257_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__mux2_1
Xhold1183 _14202_/Q vssd1 vssd1 vccd1 vccd1 hold1183/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _11850_/X vssd1 vssd1 vccd1 vccd1 _14673_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _15270_/CLK hold570/X vssd1 vssd1 vccd1 vccd1 hold569/A sky130_fd_sc_hd__dfxtp_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ hold997/X _13729_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 hold998/A sky130_fd_sc_hd__mux2_1
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _15265_/CLK hold186/X vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__dfxtp_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12884__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ hold1579/X _13512_/A0 _11779_/S vssd1 vssd1 vccd1 vccd1 _11773_/X sky130_fd_sc_hd__mux2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13512_ _13512_/A0 hold2027/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13512_/X sky130_fd_sc_hd__mux2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _10721_/X _10722_/Y _10543_/Y _10548_/C vssd1 vssd1 vccd1 vccd1 _10724_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _15426_/CLK _14492_/D vssd1 vssd1 vccd1 vccd1 _14492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13443_ _06916_/A _13450_/A _13442_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15215_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10655_ _11605_/A _11537_/A _11623_/B _15207_/Q vssd1 vssd1 vccd1 vccd1 _10656_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08382__B _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07279__A _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13593__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13374_ _13381_/A _13374_/B vssd1 vssd1 vccd1 vccd1 _15165_/D sky130_fd_sc_hd__nor2_1
XANTENNA__09261__B1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ _14356_/Q hold433/A _14420_/Q _14132_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _10587_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10946__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15113_ _15116_/CLK _15113_/D vssd1 vssd1 vccd1 vccd1 _15113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ _12330_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12354_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09239__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15044_ _15268_/CLK _15044_/D vssd1 vssd1 vccd1 vccd1 _15044_/Q sky130_fd_sc_hd__dfxtp_1
X_12256_ _12256_/A _12256_/B vssd1 vssd1 vccd1 vccd1 _12256_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06911__A _15342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _11207_/A _11207_/B _11386_/B vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_103_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10433__A _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ _12120_/A _12195_/A2 _12186_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11138_ _11320_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11138_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11963__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12546__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _10885_/B _10887_/B _11067_/X _11068_/Y vssd1 vssd1 vccd1 vccd1 _11069_/Y
+ sky130_fd_sc_hd__a211oi_2
Xclkbuf_leaf_0_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15265_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14828_ _14876_/CLK _14828_/D vssd1 vssd1 vccd1 vccd1 _14828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11426__A2 _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14759_ _15400_/CLK hold184/X vssd1 vssd1 vccd1 vccd1 _14759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07300_ _15219_/Q _11563_/B vssd1 vssd1 vccd1 vccd1 _07302_/A sky130_fd_sc_hd__or2_1
XANTENNA__09669__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ _08877_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_188_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07231_ _15201_/Q _11550_/A vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__and2_1
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__B _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07162_ _13729_/A1 hold1361/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07162_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2734_A _13428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07093_ _13729_/A1 hold2095/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07093_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11439__A _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12034__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__A2 _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07128__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ _10430_/B1 _09796_/Y _09798_/Y _09800_/Y _09802_/Y vssd1 vssd1 vccd1 vccd1
+ _09803_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ _08065_/A _07995_/B vssd1 vssd1 vccd1 vccd1 _07995_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout385_A _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _09734_/A _09734_/B _09734_/C vssd1 vssd1 vccd1 vccd1 _09734_/Y sky130_fd_sc_hd__nor3_4
XANTENNA__13103__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ _13287_/A vssd1 vssd1 vccd1 vccd1 _06946_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_179_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12862__A1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08616_ _08616_/A _08616_/B _08616_/C vssd1 vssd1 vccd1 vccd1 _08617_/C sky130_fd_sc_hd__and3_1
X_09596_ _09592_/X _09593_/Y _09451_/X _09453_/Y vssd1 vssd1 vccd1 vccd1 _09597_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ hold253/A hold817/A _14600_/Q _13969_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08547_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout817_A _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07798__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _09026_/B _08702_/B _09437_/A _08908_/A vssd1 vssd1 vccd1 vccd1 _08480_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07429_ _07429_/A _07450_/B vssd1 vssd1 vccd1 vccd1 _14059_/D sky130_fd_sc_hd__and2_1
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _11578_/A _11573_/B _14966_/Q _11580_/A vssd1 vssd1 vccd1 vccd1 _10440_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12473__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10371_ _10367_/X _10368_/Y _10191_/X _10193_/Y vssd1 vssd1 vccd1 vccd1 _10373_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _14995_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12110_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_66_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ hold885/A _14137_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08349__A2 _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _12059_/A _12041_/B vssd1 vssd1 vccd1 vccd1 _14833_/D sky130_fd_sc_hd__and2_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11353__A1 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout760 _11561_/A vssd1 vssd1 vccd1 vccd1 _11351_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__11783__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 _14946_/Q vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout782 _14943_/Q vssd1 vssd1 vccd1 vccd1 _11335_/A sky130_fd_sc_hd__buf_4
X_13992_ _15263_/CLK _13992_/D vssd1 vssd1 vccd1 vccd1 _13992_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_184_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 hold2782/X vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__buf_6
XFILLER_0_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09849__A2 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07562__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _13098_/S1 _12940_/X _12942_/X vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__a21o_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12853__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__B _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07281__B _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _13884_/Q hold675/A _13852_/Q _13820_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12874_/X sky130_fd_sc_hd__mux4_1
XANTENNA_120 _13203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_153 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613_ _15090_/CLK hold312/X vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__dfxtp_1
X_11825_ hold363/X _13679_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold364/A sky130_fd_sc_hd__mux2_1
XANTENNA__12605__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_164 _13460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_175 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13503__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10616__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_197 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14544_ _15444_/CLK _14544_/D vssd1 vssd1 vccd1 vccd1 _14544_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12700__S1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ _13742_/A1 hold983/X _11761_/S vssd1 vssd1 vccd1 vccd1 hold984/A sky130_fd_sc_hd__mux2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_79_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07501__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10707_ _10707_/A _10707_/B _10707_/C vssd1 vssd1 vccd1 vccd1 _10707_/Y sky130_fd_sc_hd__nand3_1
X_14475_ _15449_/CLK _14475_/D vssd1 vssd1 vccd1 vccd1 _14475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11687_ input46/X _13648_/B vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__or2_1
XANTENNA__10428__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_122_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13426_ _13440_/S _13426_/B vssd1 vssd1 vccd1 vccd1 _13426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ _11614_/A _10830_/B _11378_/C _11586_/A vssd1 vssd1 vccd1 vccd1 _10639_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13030__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12464__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11041__B1 _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13357_ _13360_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _15148_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10569_ _11108_/A _10746_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__o21a_1
X_12308_ _12308_/A _12308_/B _12308_/C _12308_/D vssd1 vssd1 vccd1 vccd1 _12330_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__08993__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ input135/X fanout5/X fanout3/X input103/X vssd1 vssd1 vccd1 vccd1 _13288_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_137_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15027_ _15188_/CLK _15027_/D vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13333__A2 fanout6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__B _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ _12233_/A _12236_/X _12238_/X vssd1 vssd1 vccd1 vccd1 _12239_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2609 _15115_/Q vssd1 vssd1 vccd1 vccd1 hold2609/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_leaf_17_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1908 _07508_/X vssd1 vssd1 vccd1 vccd1 _14136_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1919 _13962_/Q vssd1 vssd1 vccd1 vccd1 hold1919/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13474__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07780_ hold1091/X _13718_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 _07780_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 dmemresp_rdata[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12844__A1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09450_ _09591_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11425__C _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08401_ _08401_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_149_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09381_ _09381_/A vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__inv_2
XFILLER_0_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08332_ _08331_/B _08331_/C _08331_/A vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__10607__A1_N _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08263_ _08352_/B _08352_/C vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__and2_1
XANTENNA__10338__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07214_ hold1147/X _13715_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 _07214_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08194_ _08201_/A _08191_/X _08193_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _08195_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07145_ _13680_/A1 hold1741/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07145_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09846__B _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07076_ _13681_/A1 hold1869/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07076_/X sky130_fd_sc_hd__mux2_1
Xoutput330 _14828_/Q vssd1 vssd1 vccd1 vccd1 out2[15] sky130_fd_sc_hd__buf_12
Xoutput341 _14838_/Q vssd1 vssd1 vccd1 vccd1 out2[25] sky130_fd_sc_hd__buf_12
XFILLER_0_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12272__B _13430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput352 _14819_/Q vssd1 vssd1 vccd1 vccd1 out2[6] sky130_fd_sc_hd__buf_12
XANTENNA__12758__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09284__D _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout767_A _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13384__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _08042_/B _14426_/Q vssd1 vssd1 vccd1 vccd1 _07978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _09570_/X _09572_/X _09715_/Y _09716_/X vssd1 vssd1 vccd1 vccd1 _09717_/X
+ sky130_fd_sc_hd__o211a_1
X_06929_ _14092_/Q vssd1 vssd1 vccd1 vccd1 _06972_/B sky130_fd_sc_hd__inv_2
XANTENNA__10520__B _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _15410_/Q _14545_/Q hold933/A _14769_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09648_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07937__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ hold781/A _14117_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11351__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _11541_/A _15222_/Q vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10248__A _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _14958_/CLK hold434/X vssd1 vssd1 vccd1 vccd1 hold433/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _11281_/A _11281_/B _11280_/A _11279_/Y _11471_/B vssd1 vssd1 vccd1 vccd1
+ _11473_/C sky130_fd_sc_hd__o311ai_4
XFILLER_0_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13012__A1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12446__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11778__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ hold1021/X _13690_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__mux2_1
X_10423_ _14355_/Q hold567/A hold547/A _14131_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10424_/B sky130_fd_sc_hd__mux4_1
X_14191_ _15188_/CLK hold210/X vssd1 vssd1 vccd1 vccd1 _14191_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12997__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07557__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ _13455_/A _13142_/B vssd1 vssd1 vccd1 vccd1 _15007_/D sky130_fd_sc_hd__and2_2
X_10354_ _11541_/A _11561_/A _10830_/B _10356_/C _10185_/X vssd1 vssd1 vccd1 vccd1
+ _10362_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_21_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07276__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12749__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ hold213/A _14328_/Q hold353/A _13988_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _13073_/X sky130_fd_sc_hd__mux4_1
X_10285_ _10285_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12024_ _14985_/Q hold2672/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09772__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__A2 _08743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13079__A1 _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _09809_/C vssd1 vssd1 vccd1 vccd1 _10356_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07292__A _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__B _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13975_ _15373_/CLK _13975_/D vssd1 vssd1 vccd1 vccd1 _13975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07928__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11245__C _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ _13101_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12927_/C sky130_fd_sc_hd__or2_1
XANTENNA__12921__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ _13171_/A _12857_/B vssd1 vssd1 vccd1 vccd1 _14962_/D sky130_fd_sc_hd__nor2_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11542__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13233__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ hold1697/X _13662_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ _12917_/B1 _12783_/X _12787_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12795_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _13725_/A1 hold1785/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11739_/X sky130_fd_sc_hd__mux2_1
X_14527_ _15429_/CLK hold480/X vssd1 vssd1 vccd1 vccd1 _14527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09207__B1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _15429_/CLK _14458_/D vssd1 vssd1 vccd1 vccd1 _14458_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13003__B2 _13199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13409_ _13409_/A _13409_/B vssd1 vssd1 vccd1 vccd1 _15198_/D sky130_fd_sc_hd__and2_1
XFILLER_0_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14389_ _15385_/CLK _14389_/D vssd1 vssd1 vccd1 vccd1 _14389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07467__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08950_ _08950_/A _08997_/A _08950_/C vssd1 vssd1 vccd1 vccd1 _08997_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11317__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07901_ _07900_/B _13376_/B _12259_/A1 _13174_/B vssd1 vssd1 vccd1 vccd1 _07901_/X
+ sky130_fd_sc_hd__a22o_1
Xhold2406 hold2833/X vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__buf_1
Xhold2417 _14070_/Q vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08881_ _08866_/Y _08871_/Y _08880_/X _12241_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08882_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2428 _15313_/Q vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__buf_1
Xhold2439 _14990_/Q vssd1 vssd1 vccd1 vccd1 hold2439/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13408__S _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1705 _13999_/Q vssd1 vssd1 vccd1 vccd1 hold1705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1716 _11952_/X vssd1 vssd1 vccd1 vccd1 _14772_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07832_ _12247_/A _07832_/B vssd1 vssd1 vccd1 vccd1 _07832_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10621__A _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1727 _14119_/Q vssd1 vssd1 vccd1 vccd1 hold1727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 _11916_/X vssd1 vssd1 vccd1 vccd1 _14737_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1749 _13966_/Q vssd1 vssd1 vccd1 vccd1 hold1749/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09369__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _13668_/A1 hold1373/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07763_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12817__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09502_ _09514_/A _09501_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_78_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10828__B1 _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07694_ hold1125/X _13519_/A0 _07709_/S vssd1 vssd1 vccd1 vccd1 _07694_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09433_ _10033_/A _09864_/C _09864_/D _09435_/A vssd1 vssd1 vccd1 vccd1 _09437_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08249__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _10244_/A _09364_/B vssd1 vssd1 vccd1 vccd1 _09364_/X sky130_fd_sc_hd__or2_1
XFILLER_0_192_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12267__B _13420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ _08314_/B _08314_/C _08314_/A vssd1 vssd1 vccd1 vccd1 _08317_/D sky130_fd_sc_hd__a21o_1
XANTENNA__11171__B _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09295_ _09295_/A _09295_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_hold1198_A _13475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_42 _15205_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08246_ _10397_/A _08242_/X _08243_/X _12256_/A _06939_/Y vssd1 vssd1 vccd1 vccd1
+ _08246_/X sky130_fd_sc_hd__o32a_1
XANTENNA_53 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_64 _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_75 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11005__B1 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_86 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_97 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13379__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _08109_/A _08106_/Y _08108_/B vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__A2 _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12753__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ _13729_/A1 hold2207/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07128_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout884_A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10764__C1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07059_ _13664_/A1 hold1199/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_203_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11308__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput171 _15183_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[18] sky130_fd_sc_hd__buf_12
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput182 _15193_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[28] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ _09910_/A _10071_/A _10071_/B vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__o21bai_1
Xoutput193 _15174_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[9] sky130_fd_sc_hd__buf_12
XFILLER_0_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12600__S0 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ hold185/X vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ _10972_/A _10972_/B _10972_/C vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12711_ _12917_/A1 _12710_/X _12844_/A1 vssd1 vssd1 vccd1 vccd1 _12711_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13691_ hold519/X _13691_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 hold520/A sky130_fd_sc_hd__mux2_1
XFILLER_0_195_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ _12642_/A1 _12641_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12642_/X sky130_fd_sc_hd__a21o_1
X_15430_ _15434_/CLK _15430_/D vssd1 vssd1 vccd1 vccd1 _15430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07051__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11244__B1 _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15361_ _15361_/CLK _15361_/D vssd1 vssd1 vccd1 vccd1 _15361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12573_ hold229/A hold505/A _14599_/Q _13968_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12573_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07999__B1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10598__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _11524_/A _11524_/B vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14312_ _15367_/CLK _14312_/D vssd1 vssd1 vccd1 vccd1 _14312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12992__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15292_ _15292_/CLK hold770/X vssd1 vssd1 vccd1 vccd1 hold769/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14243_ _15436_/CLK _14243_/D vssd1 vssd1 vccd1 vccd1 _14243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11455_ _11455_/A _11455_/B vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10406_ _10406_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10746_/A sky130_fd_sc_hd__nand2_1
X_14174_ _15268_/CLK hold234/X vssd1 vssd1 vccd1 vccd1 _14174_/Q sky130_fd_sc_hd__dfxtp_1
X_11386_ _11386_/A _11386_/B vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ _13492_/A hold75/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__and2_1
X_10337_ _10380_/B vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08963__A2 _13388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _07355_/Y _13169_/B _08637_/Y vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__o21a_1
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__and2_1
XFILLER_0_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12007_ _12063_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _14816_/D sky130_fd_sc_hd__and2_1
XANTENNA__13228__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__A _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10199_ _10199_/A vssd1 vssd1 vccd1 vccd1 _10199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08271__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10798__D _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11971__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13958_ _14557_/CLK _13958_/D vssd1 vssd1 vccd1 vccd1 _13958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12909_ hold355/X _13918_/Q _12915_/S vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13889_ _15385_/CLK _13889_/D vssd1 vssd1 vccd1 vccd1 _13889_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12368__A _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12658__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ _08097_/X _08098_/Y _08099_/Y vssd1 vssd1 vccd1 vccd1 _08100_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_127_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _11288_/A1 _09079_/Y _08996_/X vssd1 vssd1 vccd1 vccd1 _12275_/B sky130_fd_sc_hd__a21o_4
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08651__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08031_ _07323_/C _08029_/X _08030_/Y vssd1 vssd1 vccd1 vccd1 _08031_/X sky130_fd_sc_hd__o21a_1
Xinput40 imemresp_data[16] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
XANTENNA__13199__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09396__B _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 imemresp_data[26] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_1
XFILLER_0_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13083__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput62 imemresp_data[7] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xhold802 hold802/A vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 in0[17] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput84 in0[27] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_1
Xhold813 hold813/A vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 in0[8] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold824 hold824/A vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 hold835/A vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold846 hold846/A vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 hold857/A vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _09982_/A _09982_/B _10182_/B vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__nand3_4
Xhold868 hold868/A vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 hold879/A vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08933_ _08933_/A vssd1 vssd1 vccd1 vccd1 _08933_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2203 _14268_/Q vssd1 vssd1 vccd1 vccd1 hold2203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2214 _07805_/X vssd1 vssd1 vccd1 vccd1 _14420_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2225 _13978_/Q vssd1 vssd1 vccd1 vccd1 hold2225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2236 _07006_/X vssd1 vssd1 vccd1 vccd1 _13825_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1502 _11744_/X vssd1 vssd1 vccd1 vccd1 _14538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2247 _14773_/Q vssd1 vssd1 vccd1 vccd1 hold2247/X sky130_fd_sc_hd__dlygate4sd3_1
X_08864_ _13876_/Q _14004_/Q _13844_/Q _13812_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08864_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10351__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1513 _14483_/Q vssd1 vssd1 vccd1 vccd1 hold1513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2258 _07150_/X vssd1 vssd1 vccd1 vccd1 _13958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2269 _14747_/Q vssd1 vssd1 vccd1 vccd1 hold2269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 _07160_/X vssd1 vssd1 vccd1 vccd1 _13968_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07136__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1535 _14390_/Q vssd1 vssd1 vccd1 vccd1 hold1535/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ _07815_/A _07815_/B vssd1 vssd1 vccd1 vccd1 _07815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11166__B _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1546 _11771_/X vssd1 vssd1 vccd1 vccd1 _14596_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ _08794_/B _08794_/C _08794_/A vssd1 vssd1 vccd1 vccd1 _08797_/B sky130_fd_sc_hd__a21o_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1557 _14640_/Q vssd1 vssd1 vccd1 vccd1 hold1557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1568 _11661_/X vssd1 vssd1 vccd1 vccd1 _14464_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_A _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1579 _14598_/Q vssd1 vssd1 vccd1 vccd1 hold1579/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07746_ _13651_/A1 hold2123/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07746_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12897__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13381__B _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07677_ _11730_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _07677_/Y sky130_fd_sc_hd__nor2_4
XANTENNA_fanout632_A _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _09413_/X _09414_/Y _09307_/X _09309_/Y vssd1 vssd1 vccd1 vccd1 _09417_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12649__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ _09347_/A _09347_/B vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _11580_/A _10010_/B _09420_/A _09277_/D vssd1 vssd1 vccd1 vccd1 _09279_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_118_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ _08312_/A _08702_/B _08228_/C _08228_/D vssd1 vssd1 vccd1 vccd1 _08230_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10526__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13074__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _11240_/A _11240_/B vssd1 vssd1 vccd1 vccd1 _11254_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _11573_/A _11594_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _11174_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ _10122_/A _10122_/B _10122_/C vssd1 vssd1 vccd1 vccd1 _10123_/D sky130_fd_sc_hd__or3_1
XANTENNA__13556__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__S _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12945__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _10056_/C vssd1 vssd1 vccd1 vccd1 _10053_/Y sky130_fd_sc_hd__inv_2
X_14930_ _15243_/CLK _14930_/D vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07046__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2770 _14492_/Q vssd1 vssd1 vccd1 vccd1 _13076_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _14973_/CLK _14861_/D vssd1 vssd1 vccd1 vccd1 _14861_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2781 _15193_/Q vssd1 vssd1 vccd1 vccd1 hold2781/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2792 _15125_/Q vssd1 vssd1 vccd1 vccd1 hold2792/X sky130_fd_sc_hd__buf_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11791__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13812_ _14731_/CLK _13812_/D vssd1 vssd1 vccd1 vccd1 _13812_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__B1 _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13454__A1 _12284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14792_ _15177_/CLK _14792_/D vssd1 vssd1 vccd1 vccd1 _14792_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07570__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09122__A2 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10955_ _10955_/A _10955_/B vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08556__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13743_ hold833/X _13743_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold834/A sky130_fd_sc_hd__mux2_1
XFILLER_0_196_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13206__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10886_ _10885_/B _10885_/C _10885_/A vssd1 vssd1 vccd1 vccd1 _10887_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_112_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13674_ hold2015/X _13674_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08881__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09505__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15413_ _15452_/CLK hold680/X vssd1 vssd1 vccd1 vccd1 hold679/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12625_ _12621_/X _12622_/X _12624_/X _12623_/X _12700_/S0 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12626_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13511__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15344_ _15424_/CLK _15344_/D vssd1 vssd1 vccd1 vccd1 _15344_/Q sky130_fd_sc_hd__dfxtp_2
X_12556_ _08435_/A _08636_/A _13149_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12557_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09976__A4 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10440__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ _11507_/A _11507_/B vssd1 vssd1 vccd1 vccd1 _11507_/X sky130_fd_sc_hd__or2_1
XANTENNA__10440__B2 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12487_ _12599_/S1 _12484_/X _12486_/X vssd1 vssd1 vccd1 vccd1 _12487_/X sky130_fd_sc_hd__a21o_1
X_15275_ _15441_/CLK _15275_/D vssd1 vssd1 vccd1 vccd1 _15275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12717__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _11598_/A _11590_/A _11573_/B _14966_/Q vssd1 vssd1 vccd1 vccd1 _11439_/D
+ sky130_fd_sc_hd__nand4_1
X_14226_ _15448_/CLK _14226_/D vssd1 vssd1 vccd1 vccd1 _14226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12193__A1 hold2610/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11966__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14157_ _15446_/CLK hold418/X vssd1 vssd1 vccd1 vccd1 hold417/A sky130_fd_sc_hd__dfxtp_1
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12651__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ _13499_/A hold63/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__and2_1
X_14088_ _15293_/CLK _14088_/D vssd1 vssd1 vccd1 vccd1 _14088_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13466__B _13466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ hold813/X _14231_/Q hold825/A _14485_/Q _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13039_/X sky130_fd_sc_hd__mux4_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09960__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07600_ _13739_/A1 hold2165/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07600_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_135_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ _08598_/B _08580_/B vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__or2_1
XFILLER_0_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09649__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10259__A1 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ hold305/X _13735_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__mux2_1
XANTENNA__08547__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__B2 _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12098__A _14989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ hold237/X _13535_/B vssd1 vssd1 vccd1 vccd1 hold238/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ _09201_/A _09201_/B vssd1 vssd1 vccd1 vccd1 _09202_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07393_ _07393_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _07393_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12826__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09132_ _10126_/A _09131_/X _09130_/X vssd1 vssd1 vccd1 vccd1 _09133_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12956__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10431__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ _09060_/Y _09061_/X _08944_/B _08944_/Y vssd1 vssd1 vccd1 vccd1 _09064_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10346__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08014_ _08014_/A _08014_/B _08014_/C vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold610 hold610/A vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 hold621/A vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08388__B1 _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 hold632/A vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08927__A2 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold643 hold643/A vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold654 hold654/A vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold665 hold665/A vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 hold676/A vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold687 hold687/A vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 hold698/A vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13376__B _13376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09965_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout582_A _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2000 _07030_/X vssd1 vssd1 vccd1 vccd1 _13847_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12280__B _13446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2011 _15265_/Q vssd1 vssd1 vccd1 vccd1 hold2011/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2022 _07026_/X vssd1 vssd1 vccd1 vccd1 _13843_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08916_ _08917_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _08916_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10081__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2033 _15438_/Q vssd1 vssd1 vccd1 vccd1 hold2033/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2044 _07501_/X vssd1 vssd1 vccd1 vccd1 _14129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09896_ _09896_/A _09896_/B _09896_/C _09896_/D vssd1 vssd1 vccd1 vccd1 _09896_/Y
+ sky130_fd_sc_hd__nor4_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2055 _14035_/Q vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _11932_/X vssd1 vssd1 vccd1 vccd1 _14752_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _15282_/Q vssd1 vssd1 vccd1 vccd1 hold1321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2066 _11819_/X vssd1 vssd1 vccd1 vccd1 _14643_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2077 _14066_/Q vssd1 vssd1 vccd1 vccd1 _07408_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 _13680_/X vssd1 vssd1 vccd1 vccd1 _15387_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ _12221_/B _08845_/X _08846_/Y _08844_/X vssd1 vssd1 vccd1 vccd1 _13387_/B
+ sky130_fd_sc_hd__a31o_4
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2088 _11908_/X vssd1 vssd1 vccd1 vccd1 _14729_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _13957_/Q vssd1 vssd1 vccd1 vccd1 hold1343/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07363__A1 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1354 _11901_/X vssd1 vssd1 vccd1 vccd1 _14722_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout847_A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2099 _14502_/Q vssd1 vssd1 vccd1 vccd1 hold2099/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13392__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1365 _15385_/Q vssd1 vssd1 vccd1 vccd1 hold1365/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1376 _11707_/X vssd1 vssd1 vccd1 vccd1 _14503_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ _08778_/A _08778_/B vssd1 vssd1 vccd1 vccd1 _08788_/A sky130_fd_sc_hd__xor2_2
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1387 _13882_/Q vssd1 vssd1 vccd1 vccd1 hold1387/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13436__A1 _12275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _11781_/X vssd1 vssd1 vccd1 vccd1 _14606_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__A _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ hold1619/X _13735_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07729_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12644__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10740_ _10951_/B _10599_/X _10601_/X _11640_/B1 vssd1 vssd1 vccd1 vccd1 _10740_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ _10496_/A _10498_/B _10669_/A _10670_/Y vssd1 vssd1 vccd1 vccd1 _10673_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12410_ _14657_/Q _13930_/Q _12459_/S vssd1 vssd1 vccd1 vccd1 _12410_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13390_ _13390_/A _13390_/B vssd1 vssd1 vccd1 vccd1 _15181_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ _12366_/A _12341_/B vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__or2_1
XFILLER_0_180_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13047__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ _15377_/CLK _15060_/D vssd1 vssd1 vccd1 vccd1 _15060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12272_ _13150_/A _13430_/B vssd1 vssd1 vccd1 vccd1 _14921_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08379__B1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ _15379_/CLK hold622/X vssd1 vssd1 vccd1 vccd1 hold621/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12175__A1 hold2605/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ _11455_/B _11221_/Y _11033_/A _11035_/A vssd1 vssd1 vccd1 vccd1 _11264_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07565__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _11590_/A _11594_/B _11155_/C _11435_/A vssd1 vssd1 vccd1 vccd1 _11156_/B
+ sky130_fd_sc_hd__a22o_1
X_10105_ _11320_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10105_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07284__B _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11085_ _10900_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11087_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12478__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ _10036_/A _10036_/B _10141_/B vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__nand3_1
X_14913_ _15391_/CLK _14913_/D vssd1 vssd1 vccd1 vccd1 _14913_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09343__A2 _09342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13506__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14844_ _14844_/CLK _14844_/D vssd1 vssd1 vccd1 vccd1 _14844_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12410__S _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07504__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14775_ _14775_/CLK _14775_/D vssd1 vssd1 vccd1 vccd1 _14775_/Q sky130_fd_sc_hd__dfxtp_1
X_11987_ hold299/X _15062_/Q _11993_/S vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__mux2_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ hold1269/X _15046_/Q _13732_/S vssd1 vssd1 vccd1 vccd1 _13726_/X sky130_fd_sc_hd__mux2_1
X_10938_ _14358_/Q hold667/A _14422_/Q _14134_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _10939_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10869_ _11340_/A _15223_/Q vssd1 vssd1 vccd1 vccd1 _10870_/B sky130_fd_sc_hd__nand2_1
X_13657_ hold1023/X _13657_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 _13657_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08843__B _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11550__A _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ hold803/A _14537_/Q _14697_/Q _14761_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12608_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_183_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13588_ _13588_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__or2_1
XFILLER_0_14_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15327_ _15422_/CLK _15327_/D vssd1 vssd1 vccd1 vccd1 _15327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10166__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ hold1161/X hold577/X hold2808/X hold2109/X _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12539_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15258_ _15258_/CLK _15258_/D vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ _15040_/CLK hold802/X vssd1 vssd1 vccd1 vccd1 hold801/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13477__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15189_ _15190_/CLK _15189_/D vssd1 vssd1 vccd1 vccd1 _15189_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13196__B _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _07149_/X vssd1 vssd1 vccd1 vccd1 _07181_/S sky130_fd_sc_hd__clkbuf_16
Xfanout419 _13650_/Y vssd1 vssd1 vccd1 vccd1 _13666_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _09747_/X _09748_/Y _09557_/X _09602_/A vssd1 vssd1 vccd1 vccd1 _09750_/X
+ sky130_fd_sc_hd__a211o_1
X_06962_ hold237/A hold273/A _06962_/C _06961_/X vssd1 vssd1 vccd1 vccd1 _06962_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__11126__C1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _10033_/A _08809_/B _08809_/D _09138_/A vssd1 vssd1 vccd1 vccd1 _08703_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11677__A0 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _09681_/A _09681_/B _09681_/C vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08632_ _08526_/B _08630_/Y _08631_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _08632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08563_ _08981_/A _08562_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _08563_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09098__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07514_ hold1003/X hold2816/X _07528_/S vssd1 vssd1 vccd1 vccd1 _07514_/X sky130_fd_sc_hd__mux2_1
X_08494_ _08776_/B _08809_/B _08809_/D _08776_/A vssd1 vssd1 vccd1 vccd1 _08496_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07445_ _08345_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _14075_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout428_A _11829_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08058__C1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ _06909_/Y _14062_/Q _07405_/A _15345_/Q vssd1 vssd1 vccd1 vccd1 _07376_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12275__B _12275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09115_ hold2747/X input8/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ _09167_/B _09045_/C _09045_/A vssd1 vssd1 vccd1 vccd1 _09047_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09865__A _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__C _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12157__A1 _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout797_A _14490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13387__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14921__D _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 hold440/A vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__A _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold451 hold451/A vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 hold462/A vssd1 vssd1 vccd1 vccd1 hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold473/A vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold484 hold484/A vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/A vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13106__B1 _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ hold445/A _13948_/Q _15449_/Q _13916_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _09949_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _09879_/A _09879_/B _10030_/B vssd1 vssd1 vccd1 vccd1 _09881_/B sky130_fd_sc_hd__nand3_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 _07041_/X vssd1 vssd1 vccd1 vccd1 _13858_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 _14634_/Q vssd1 vssd1 vccd1 vccd1 hold1151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _13665_/A1 hold1635/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__mux2_1
Xhold1162 _07654_/X vssd1 vssd1 vccd1 vccd1 _14275_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1173 _14769_/Q vssd1 vssd1 vccd1 vccd1 hold1173/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12230__S _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ hold841/A _14129_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12890_/X sky130_fd_sc_hd__mux2_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 _07578_/X vssd1 vssd1 vccd1 vccd1 _14202_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 _14601_/Q vssd1 vssd1 vccd1 vccd1 hold1195/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ hold1249/X _13728_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__mux2_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _15072_/CLK hold204/X vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__dfxtp_1
X_11772_ hold1317/X _13725_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_138_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10543_/Y _10548_/C _10721_/X _10722_/Y vssd1 vssd1 vccd1 vccd1 _10723_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13659_/A1 hold1417/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13511_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _15324_/CLK _14491_/D vssd1 vssd1 vccd1 vccd1 _14491_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ _11569_/A _11605_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _10836_/A
+ sky130_fd_sc_hd__nand4_1
X_13442_ _13450_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13442_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__B _14965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ _13373_/A _13373_/B _13373_/C vssd1 vssd1 vccd1 vccd1 _15164_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_181_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09261__A1 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ _11509_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09261__B2 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15112_ _15116_/CLK _15112_/D vssd1 vssd1 vccd1 vccd1 _15112_/Q sky130_fd_sc_hd__dfxtp_1
X_12324_ _12325_/B vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__inv_2
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12255_ _10873_/A _08892_/A _08312_/A _08677_/A vssd1 vssd1 vccd1 vccd1 _12256_/B
+ sky130_fd_sc_hd__a22o_1
X_15043_ _15433_/CLK _15043_/D vssd1 vssd1 vccd1 vccd1 hold465/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08447__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07295__A _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _11390_/A _11623_/A _11206_/C _11386_/A vssd1 vssd1 vccd1 vccd1 _11386_/B
+ sky130_fd_sc_hd__nand4_1
X_12186_ _14904_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__or2_1
XANTENNA_output347_A _14843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11137_ _11122_/Y _11127_/Y _11136_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _11138_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11068_ _11240_/B _11067_/C _11067_/A vssd1 vssd1 vccd1 vccd1 _11068_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13236__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _10129_/A _10827_/C _10019_/C _10019_/D vssd1 vssd1 vccd1 vccd1 _10020_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_188_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14827_ _14844_/CLK _14827_/D vssd1 vssd1 vccd1 vccd1 _14827_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10882__A1 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11506__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14758_ _15045_/CLK _14758_/D vssd1 vssd1 vccd1 vccd1 _14758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ hold419/X _13742_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold420/A sky130_fd_sc_hd__mux2_1
XFILLER_0_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09669__B _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14689_ _15394_/CLK hold672/X vssd1 vssd1 vccd1 vccd1 hold671/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07230_ _07230_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__and2_1
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12387__A1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08292__C _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07161_ _13662_/A1 hold1899/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10398__B1 _11474_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ _13728_/A1 hold2273/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07092_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12139__A1 hold2586/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2727_A _15187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11439__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09802_ _10244_/A _09801_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09802_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13639__A1 _08179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07994_ _14270_/Q _14206_/Q hold751/A _14460_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07995_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_199_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09733_ _09733_/A _09733_/B _09733_/C vssd1 vssd1 vccd1 vccd1 _09734_/C sky130_fd_sc_hd__nor3_2
X_06945_ _14094_/Q vssd1 vssd1 vccd1 vccd1 _12128_/B sky130_fd_sc_hd__inv_2
XFILLER_0_207_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12050__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _09663_/A _09813_/B _09663_/C vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ _08616_/A _08616_/B _08616_/C vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09595_ _09451_/X _09453_/Y _09592_/X _09593_/Y vssd1 vssd1 vccd1 vccd1 _09597_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout545_A _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06983__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ _08856_/C _08545_/Y _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08546_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08764__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08477_ _09661_/A _08685_/C vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__and2_1
XANTENNA_fanout712_A _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ _07428_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _14058_/D sky130_fd_sc_hd__and2_1
XFILLER_0_163_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07359_ _07359_/A _07359_/B _07910_/B _07358_/X vssd1 vssd1 vccd1 vccd1 _07359_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_163_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12473__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ _10373_/B vssd1 vssd1 vccd1 vccd1 _10370_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ _08909_/A _08909_/B _08909_/C vssd1 vssd1 vccd1 vccd1 _09030_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12040_ hold2591/X hold2690/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A2 _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 _14952_/Q vssd1 vssd1 vccd1 vccd1 _10306_/A sky130_fd_sc_hd__buf_2
Xfanout761 _08809_/D vssd1 vssd1 vccd1 vccd1 _09979_/B sky130_fd_sc_hd__buf_6
Xfanout772 _11333_/B vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13564__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout783 _11340_/A vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__buf_4
XANTENNA__12838__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13991_ _15427_/CLK _13991_/D vssd1 vssd1 vccd1 vccd1 _13991_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout794 _12988_/C1 vssd1 vssd1 vccd1 vccd1 _06944_/A sky130_fd_sc_hd__buf_8
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12942_ _13092_/A1 _12941_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_176_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12853__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07054__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _15209_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ hold205/A hold559/A hold507/A _13980_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12873_/X sky130_fd_sc_hd__mux4_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _13144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14612_ _14612_/CLK _14612_/D vssd1 vssd1 vccd1 vccd1 _14612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11824_ hold481/X _13711_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold482/A sky130_fd_sc_hd__mux2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _13437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_176 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10616__A1 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_187 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10616__B2 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_198 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ _15377_/CLK _14543_/D vssd1 vssd1 vccd1 vccd1 _14543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _13708_/A1 hold1149/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11755_/X sky130_fd_sc_hd__mux2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ _10707_/A _10707_/B _10707_/C vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__and3_1
XFILLER_0_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14474_ _15445_/CLK hold588/X vssd1 vssd1 vccd1 vccd1 hold587/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _06907_/A _11650_/B _11685_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _14488_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13425_ _08435_/B _13450_/A _13424_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _13425_/X
+ sky130_fd_sc_hd__o211a_1
X_10637_ _11586_/A _11614_/A _10830_/B _11378_/C vssd1 vssd1 vccd1 vccd1 _10639_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12464__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10919__A2 _10918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11041__A1 _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__B2 _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08442__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13356_ _13360_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _15147_/D sky130_fd_sc_hd__nor2_1
X_10568_ _10744_/A _10568_/B vssd1 vssd1 vccd1 vccd1 _10746_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _15349_/Q _06937_/Y _07841_/X _12306_/X vssd1 vssd1 vccd1 vccd1 _12308_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13287_ _13287_/A _13287_/B vssd1 vssd1 vccd1 vccd1 _15115_/D sky130_fd_sc_hd__nor2_1
X_10499_ _10498_/B _10498_/C _10498_/A vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__o21ai_2
X_15026_ _15188_/CLK _15026_/D vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__dfxtp_1
X_12238_ _12231_/A _12237_/X _12243_/A vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11974__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__C1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12102_/A _12173_/A2 _12168_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1909 _14609_/Q vssd1 vssd1 vccd1 vccd1 hold1909/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_127_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 dmemresp_rdata[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07472__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11425__D _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08400_ _09164_/A _09712_/A _08468_/A _08400_/D vssd1 vssd1 vccd1 vccd1 _08468_/B
+ sky130_fd_sc_hd__nand4_2
X_09380_ _10351_/A _09809_/C _09295_/A _09292_/X vssd1 vssd1 vccd1 vccd1 _09381_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08331_ _08331_/A _08331_/B _08331_/C vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_129_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10619__A _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08262_ _08257_/A _08441_/B _08250_/Y _08261_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1
+ _08262_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_184_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10338__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07213_ hold401/X _13681_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold402/A sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08193_ _08197_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08193_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08659__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07144_ _13745_/A1 hold1957/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07144_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09846__C _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12780__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ _13680_/A1 hold1913/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07075_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput320 _14851_/Q vssd1 vssd1 vccd1 vccd1 out1[6] sky130_fd_sc_hd__buf_12
Xoutput331 _14829_/Q vssd1 vssd1 vccd1 vccd1 out2[16] sky130_fd_sc_hd__buf_12
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput342 _14839_/Q vssd1 vssd1 vccd1 vccd1 out2[26] sky130_fd_sc_hd__buf_12
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07139__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput353 _14820_/Q vssd1 vssd1 vccd1 vccd1 out2[7] sky130_fd_sc_hd__buf_12
XANTENNA__11884__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13384__B _13384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__C _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _13750_/A _13345_/B vssd1 vssd1 vccd1 vccd1 _07981_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_199_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09716_ _09715_/B _09715_/C _09715_/A vssd1 vssd1 vccd1 vccd1 _09716_/X sky130_fd_sc_hd__a21o_1
X_06928_ _14082_/Q vssd1 vssd1 vccd1 vccd1 _06928_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09647_ _10426_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09647_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12048__A0 _12114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07602__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__C _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08529_ _08530_/A _08530_/C _08530_/D _08530_/B vssd1 vssd1 vccd1 vccd1 _08569_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_195_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11351__C _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _11540_/A _11540_/B vssd1 vssd1 vccd1 vccd1 _11548_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout5_A fanout6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11473_/B sky130_fd_sc_hd__or2_1
XFILLER_0_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12446__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12220__A0 hold2757/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ hold1473/X _13656_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__mux2_1
X_10422_ _11509_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10422_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_122_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14190_ _15188_/CLK hold182/X vssd1 vssd1 vccd1 vccd1 _14190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10353_ _10140_/A _10139_/B _10137_/X vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__a21o_1
X_13141_ _13381_/A _13141_/B vssd1 vssd1 vccd1 vccd1 _15006_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07049__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ _14811_/Q hold875/A hold341/A _14747_/Q _13066_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _13072_/X sky130_fd_sc_hd__mux4_1
X_10284_ _11590_/A _10283_/C _11570_/B _11598_/A vssd1 vssd1 vccd1 vccd1 _10285_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ _12059_/A _12023_/B vssd1 vssd1 vccd1 vccd1 _14824_/D sky130_fd_sc_hd__and2_1
XANTENNA__11794__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__C1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07573__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13079__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout580 _15219_/Q vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__buf_6
XFILLER_0_75_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07292__B _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout591 _15214_/Q vssd1 vssd1 vccd1 vccd1 _09809_/C sky130_fd_sc_hd__buf_4
X_13974_ _15375_/CLK _13974_/D vssd1 vssd1 vccd1 vccd1 _13974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09152__B1 _15210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ _12921_/X _12922_/X _12924_/X _12923_/X _12950_/S0 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12926_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11245__D _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _13106_/A1 _13161_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12857_/B sky130_fd_sc_hd__o21a_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11542__B _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ hold1057/X _13661_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11807_/X sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12899_/S1 _12784_/X _12786_/X vssd1 vssd1 vccd1 vccd1 _12787_/X sky130_fd_sc_hd__a21o_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14750_/CLK _14526_/D vssd1 vssd1 vccd1 vccd1 _14526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11738_ _13691_/A1 hold901/X _11745_/S vssd1 vssd1 vccd1 vccd1 hold902/A sky130_fd_sc_hd__mux2_1
XFILLER_0_138_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11969__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09207__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ _15360_/CLK _14457_/D vssd1 vssd1 vccd1 vccd1 _14457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11669_ _13700_/A1 hold1623/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13003__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08851__B _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13408_ _07908_/A _12261_/B _13468_/A vssd1 vssd1 vccd1 vccd1 _13409_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14388_ _15453_/CLK _14388_/D vssd1 vssd1 vccd1 vccd1 _14388_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12762__A1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13339_ _08637_/B _07912_/X hold2354/X vssd1 vssd1 vccd1 vccd1 _13339_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__B1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15009_ _15268_/CLK _15009_/D vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__dfxtp_1
X_07900_ _07900_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _07900_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_110_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2407 _13561_/X vssd1 vssd1 vccd1 vccd1 _15306_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2418 _14859_/Q vssd1 vssd1 vccd1 vccd1 hold2418/X sky130_fd_sc_hd__dlygate4sd3_1
X_08880_ _08880_/A1 _08873_/Y _08875_/Y _08877_/Y _08879_/Y vssd1 vssd1 vccd1 vccd1
+ _08880_/X sky130_fd_sc_hd__o32a_1
XANTENNA__08194__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2429 _13575_/X vssd1 vssd1 vccd1 vccd1 _15313_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1706 _07192_/X vssd1 vssd1 vccd1 vccd1 _13999_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07831_ hold453/A hold975/A hold635/A _13896_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _07832_/B sky130_fd_sc_hd__mux4_1
Xhold1717 _13927_/Q vssd1 vssd1 vccd1 vccd1 hold1717/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10621__B _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1728 _07491_/X vssd1 vssd1 vccd1 vccd1 _14119_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _14205_/Q vssd1 vssd1 vccd1 vccd1 hold1739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07762_ _13519_/A0 hold2051/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07762_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09369__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09501_ _13881_/Q _14009_/Q hold565/A _13817_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09501_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10828__A1 _14954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2794_A _15066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10828__B2 _14953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07693_ hold1449/X _13666_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 _07693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _09432_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09203__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09363_ _14799_/Q _14511_/Q _14639_/Q _14735_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09364_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09446__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ _08314_/A _08314_/B _08314_/C vssd1 vssd1 vccd1 vccd1 _08317_/C sky130_fd_sc_hd__nand3_2
X_09294_ _10351_/A _09809_/C vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11171__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_10 _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_21 _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _08244_/A _08244_/C _08244_/B vssd1 vssd1 vccd1 vccd1 _08245_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11879__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_43 _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_54 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A _07115_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_65 clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__A1 _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_87 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11005__B2 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_183_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_98 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _07900_/B _08175_/Y _08136_/X vssd1 vssd1 vccd1 vccd1 _08176_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13379__B _13379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12283__B _13452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A2 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07127_ _13728_/A1 hold2277/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_63_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _13663_/A1 hold2179/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07058_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout877_A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13395__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 _15184_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[19] sky130_fd_sc_hd__buf_12
Xoutput183 _15194_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[29] sky130_fd_sc_hd__buf_12
XANTENNA__08489__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput194 _06951_/X vssd1 vssd1 vccd1 vccd1 dmemreq_type sky130_fd_sc_hd__buf_12
XANTENNA__12600__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_121_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12364__S0 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10970_/B _11150_/B _10970_/A vssd1 vssd1 vccd1 vccd1 _10972_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12710_ _14669_/Q _13942_/Q _12741_/S vssd1 vssd1 vccd1 vccd1 _12710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13690_ hold641/X _13690_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 hold642/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_136_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ hold989/A _14247_/Q _12641_/S vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_167_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11244__A1 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15360_ _15360_/CLK _15360_/D vssd1 vssd1 vccd1 vccd1 _15360_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_16_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__B2 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _14791_/Q _14503_/Q _14631_/Q hold967/A _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12572_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07999__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ _14602_/CLK _14311_/D vssd1 vssd1 vccd1 vccd1 _14311_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11789__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12992__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15291_ _15457_/CLK hold678/X vssd1 vssd1 vccd1 vccd1 hold677/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14242_ _14955_/CLK hold734/X vssd1 vssd1 vccd1 vccd1 hold733/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07568__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11454_ _11454_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12744__A1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _10744_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__xor2_1
X_14173_ _15268_/CLK hold212/X vssd1 vssd1 vccd1 vccd1 _14173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ _13129_/A hold25/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__and2_1
X_10336_ _10336_/A _10336_/B _10336_/C vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__and3_1
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output162_A _15165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13509__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _10267_/A _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__nor3_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13080_/A1 _13054_/X _13052_/X vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08970__A2_N _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ hold2586/X hold2668/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07507__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11537__B _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ _10198_/A _10198_/B _10198_/C vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__nor3_2
XANTENNA__08271__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13457__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13957_ _15458_/CLK _13957_/D vssd1 vssd1 vccd1 vccd1 _13957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12908_ hold2800/X _14549_/Q _14709_/Q _14773_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12908_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_158_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ _14791_/CLK _13888_/D vssd1 vssd1 vccd1 vccd1 _13888_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09023__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12839_ hold979/X _14223_/Q hold389/X hold1777/X _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12839_/X sky130_fd_sc_hd__mux4_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12658__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11699__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ _15190_/CLK _14509_/D vssd1 vssd1 vccd1 vccd1 _14509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold2375_A _15035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08030_ _07323_/C _08029_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _08030_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput30 dmemresp_rdata[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13199__B _13199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput41 imemresp_data[17] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput52 imemresp_data[27] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 imemresp_data[8] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13083__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold803 hold803/A vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold2542_A _15002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput74 in0[18] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_1
Xhold814 hold814/A vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 in0[28] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_1
Xhold825 hold825/A vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput96 in0[9] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 hold836/A vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold847 hold847/A vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 hold858/A vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _10185_/A _11378_/C _09981_/C _10182_/A vssd1 vssd1 vccd1 vccd1 _10182_/B
+ sky130_fd_sc_hd__nand4_2
Xhold869 hold869/A vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
X_08932_ _08932_/A _08932_/B _08932_/C vssd1 vssd1 vccd1 vccd1 _08933_/A sky130_fd_sc_hd__and3_2
XFILLER_0_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2204 _07647_/X vssd1 vssd1 vccd1 vccd1 _14268_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_62_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2215 _14762_/Q vssd1 vssd1 vccd1 vccd1 hold2215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2226 _07170_/X vssd1 vssd1 vccd1 vccd1 _13978_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2237 _14811_/Q vssd1 vssd1 vccd1 vccd1 hold2237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1503 _14015_/Q vssd1 vssd1 vccd1 vccd1 hold1503/X sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ hold231/A _14312_/Q _14603_/Q _13972_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08863_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10351__B _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2248 _11953_/X vssd1 vssd1 vccd1 vccd1 _14773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2259 _14467_/Q vssd1 vssd1 vccd1 vccd1 hold2259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1514 _11680_/X vssd1 vssd1 vccd1 vccd1 _14483_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 _13961_/Q vssd1 vssd1 vccd1 vccd1 hold1525/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1536 _07774_/X vssd1 vssd1 vccd1 vccd1 _14390_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07814_ hold859/A _13800_/Q _07816_/S vssd1 vssd1 vccd1 vccd1 _07815_/B sky130_fd_sc_hd__mux2_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11166__C _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1547 _13960_/Q vssd1 vssd1 vccd1 vccd1 hold1547/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08794_ _08794_/A _08794_/B _08794_/C vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__nand3_1
Xhold1558 _11816_/X vssd1 vssd1 vccd1 vccd1 _14640_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09116__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1569 _13844_/Q vssd1 vssd1 vccd1 vccd1 hold1569/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12346__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ _11652_/A _13502_/B vssd1 vssd1 vccd1 vccd1 _07745_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__12897__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A1 hold2441/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ hold1995/X _13715_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 _07676_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12278__B _13442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _09307_/X _09309_/Y _09413_/X _09414_/Y vssd1 vssd1 vccd1 vccd1 _09417_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout625_A _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12649__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06991__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _09346_/A _09346_/B _09346_/C vssd1 vssd1 vccd1 vccd1 _09347_/B sky130_fd_sc_hd__or3_1
XFILLER_0_192_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13620__C1 _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _10000_/A _10010_/B _09420_/A _09277_/D vssd1 vssd1 vccd1 vccd1 _09459_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__A _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08312_/A _08702_/B _08228_/C _08228_/D vssd1 vssd1 vccd1 vccd1 _08230_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_132_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10526__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13074__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ _08289_/A _08159_/B _08093_/A vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12821__S1 _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _11594_/A _11569_/B _11563_/B _11573_/A vssd1 vssd1 vccd1 vccd1 _11174_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10121_ _10122_/A _10122_/B _10122_/C vssd1 vssd1 vccd1 vccd1 _10328_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _10052_/A _10164_/A _10052_/C vssd1 vssd1 vccd1 vccd1 _10056_/C sky130_fd_sc_hd__nand3_2
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08012__A _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2760 _15191_/Q vssd1 vssd1 vccd1 vccd1 hold2760/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _14973_/CLK _14860_/D vssd1 vssd1 vccd1 vccd1 _14860_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2771 _13077_/X vssd1 vssd1 vccd1 vccd1 hold2771/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2782 _14492_/Q vssd1 vssd1 vccd1 vccd1 hold2782/X sky130_fd_sc_hd__buf_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2793 _15114_/Q vssd1 vssd1 vccd1 vccd1 _08843_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12337__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _15369_/CLK _13811_/D vssd1 vssd1 vccd1 vccd1 _13811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13572__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ _14791_/CLK _14791_/D vssd1 vssd1 vccd1 vccd1 _14791_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11373__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ hold437/X _13742_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold438/A sky130_fd_sc_hd__mux2_1
X_10954_ _07253_/Y _07296_/B _10599_/X _10952_/B _07255_/B vssd1 vssd1 vccd1 vccd1
+ _10955_/B sky130_fd_sc_hd__o221a_1
XANTENNA__07062__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13673_ hold551/X _13673_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold552/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10885_ _10885_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10887_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15412_ _15449_/CLK _15412_/D vssd1 vssd1 vccd1 vccd1 _15412_/Q sky130_fd_sc_hd__dfxtp_1
X_12624_ _13874_/Q hold303/A _13842_/Q _13810_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12624_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09505__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08682__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11312__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15343_ _15424_/CLK _15343_/D vssd1 vssd1 vccd1 vccd1 _15343_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12555_ _12327_/A _12554_/X _12552_/X vssd1 vssd1 vccd1 vccd1 _13149_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07298__A _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11506_ hold369/A hold385/A hold787/A hold991/A _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11507_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10440__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15274_ _15371_/CLK _15274_/D vssd1 vssd1 vccd1 vccd1 _15274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12486_ _12642_/A1 _12485_/X _12644_/A1 vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12717__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ _15062_/CLK _14225_/D vssd1 vssd1 vccd1 vccd1 _14225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _11590_/A _11573_/B _14966_/Q _11598_/A vssd1 vssd1 vccd1 vccd1 _11439_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14156_ _15445_/CLK hold306/X vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__dfxtp_1
X_11368_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13107_ _13107_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _14972_/D sky130_fd_sc_hd__nor2_1
X_10319_ _10483_/B _10318_/C _10318_/A vssd1 vssd1 vccd1 vccd1 _10320_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14087_ _15214_/CLK _14087_/D vssd1 vssd1 vccd1 vccd1 _14087_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _13750_/A _13371_/B _11298_/X vssd1 vssd1 vccd1 vccd1 _11299_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12556__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _06943_/A _13033_/X _13037_/X hold2774/X vssd1 vssd1 vccd1 vccd1 _13045_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11982__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09960__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__A _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09649__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14989_ _14989_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 _14989_/Q sky130_fd_sc_hd__dfxtp_1
X_07530_ hold2805/X hold169/X _07544_/S vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__mux2_1
XANTENNA__10259__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12653__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07461_ _07461_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07461_/X sky130_fd_sc_hd__and2_1
XFILLER_0_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_182_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15361_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09200_ _09201_/A _09201_/B vssd1 vssd1 vccd1 vccd1 _09202_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13702__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07392_ _13369_/A _07926_/A vssd1 vssd1 vccd1 vccd1 _14022_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07700__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09131_ _09571_/A _09714_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__and3_1
XANTENNA__12500__S0 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2757_A _15101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _08944_/B _08944_/Y _09060_/Y _09061_/X vssd1 vssd1 vccd1 vccd1 _09196_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10346__B _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08013_ _08312_/A _08012_/B _08012_/C _08012_/D vssd1 vssd1 vccd1 vccd1 _08014_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold600 hold600/A vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 hold611/A vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08388__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold622 hold622/A vssd1 vssd1 vccd1 vccd1 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08388__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold633 hold633/A vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07936__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold644 hold644/A vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold655 hold655/A vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 hold666/A vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold677 hold677/A vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold688/A vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__or2_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold699 hold699/A vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2001 _13977_/Q vssd1 vssd1 vccd1 vccd1 hold2001/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2012 _13507_/X vssd1 vssd1 vccd1 vccd1 _15265_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07147__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08915_ _08915_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08917_/B sky130_fd_sc_hd__xnor2_2
Xhold2023 _14500_/Q vssd1 vssd1 vccd1 vccd1 hold2023/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09895_ _10052_/A _09894_/B _09741_/A vssd1 vssd1 vccd1 vccd1 _09896_/D sky130_fd_sc_hd__o21ba_1
XANTENNA__10081__B _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2034 _13728_/X vssd1 vssd1 vccd1 vccd1 _15438_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 _07138_/X vssd1 vssd1 vccd1 vccd1 _13948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2045 _13860_/Q vssd1 vssd1 vccd1 vccd1 hold2045/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11892__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2056 _06938_/Y vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 _14291_/Q vssd1 vssd1 vccd1 vccd1 hold1311/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1322 _13524_/X vssd1 vssd1 vccd1 vccd1 _15282_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ _07323_/B _08846_/B _08846_/C vssd1 vssd1 vccd1 vccd1 _08846_/Y sky130_fd_sc_hd__nand3b_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2067 _14494_/Q vssd1 vssd1 vccd1 vccd1 hold2067/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2078 _07408_/X vssd1 vssd1 vccd1 vccd1 _14038_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06986__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1333 _15393_/Q vssd1 vssd1 vccd1 vccd1 hold1333/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12892__B1 _14490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2089 _13947_/Q vssd1 vssd1 vccd1 vccd1 hold2089/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 _07147_/X vssd1 vssd1 vccd1 vccd1 _13957_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1355 _15262_/Q vssd1 vssd1 vccd1 vccd1 hold1355/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12319__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13392__B _13392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1366 _13678_/X vssd1 vssd1 vccd1 vccd1 _15385_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1377 _14793_/Q vssd1 vssd1 vccd1 vccd1 hold1377/X sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ _14950_/Q _08776_/X _08775_/X vssd1 vssd1 vccd1 vccd1 _08778_/B sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout742_A _14954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14919__D _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1388 _07066_/X vssd1 vssd1 vccd1 vccd1 _13882_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 _14721_/Q vssd1 vssd1 vccd1 vccd1 hold1399/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ hold1675/X _13734_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07728_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_173_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15369_/CLK sky130_fd_sc_hd__clkbuf_16
X_07659_ hold799/X _13698_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold800/A sky130_fd_sc_hd__mux2_1
XFILLER_0_193_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10670_ _10668_/A _10668_/B _10464_/B vssd1 vssd1 vccd1 vccd1 _10670_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12322__B1_N _12294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09328_/B _09328_/C _09328_/A vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_153_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08076__B1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12340_ hold251/A hold743/A hold907/A _13959_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12341_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__B1 _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13047__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ _13150_/A _12271_/B vssd1 vssd1 vccd1 vccd1 _14920_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12752__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14010_ _15089_/CLK hold618/X vssd1 vssd1 vccd1 vccd1 hold617/A sky130_fd_sc_hd__dfxtp_1
X_11222_ _11033_/A _11035_/A _11455_/B _11221_/Y vssd1 vssd1 vccd1 vccd1 _11460_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__09040__A2 _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13059__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _11597_/A _11598_/A _11573_/B _14966_/Q vssd1 vssd1 vccd1 vccd1 _11435_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__10272__A _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07057__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ _10089_/Y _10094_/Y _10103_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _10105_/B sky130_fd_sc_hd__a221o_1
XANTENNA__12558__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ _11086_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11087_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11135__B1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _10142_/B _10316_/B _10035_/C _10141_/A vssd1 vssd1 vccd1 vccd1 _10141_/B
+ sky130_fd_sc_hd__nand4_1
X_14912_ _15395_/CLK _14912_/D vssd1 vssd1 vccd1 vccd1 _14912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2590 _12270_/B vssd1 vssd1 vccd1 vccd1 _13426_/B sky130_fd_sc_hd__buf_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ _14844_/CLK _14843_/D vssd1 vssd1 vccd1 vccd1 _14843_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14774_ _15452_/CLK _14774_/D vssd1 vssd1 vccd1 vccd1 _14774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ hold1857/X _13741_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__mux2_1
X_13725_ hold1543/X _13725_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__mux2_1
X_10937_ _11509_/A _10937_/B vssd1 vssd1 vccd1 vccd1 _10937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_196_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09004__C _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_164_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15442_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12927__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13522__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ hold893/X _13656_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold894/A sky130_fd_sc_hd__mux2_1
X_10868_ _10868_/A _10868_/B vssd1 vssd1 vccd1 vccd1 _10870_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06925__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07520__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12938__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09301__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11550__B _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ _12607_/A _12607_/B vssd1 vssd1 vccd1 vccd1 _14952_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08067__B1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10447__A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__A1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _10568_/B _13586_/B _13586_/Y _13409_/A vssd1 vssd1 vccd1 vccd1 _15319_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _11569_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _10801_/C sky130_fd_sc_hd__and2_1
XFILLER_0_121_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _15422_/CLK _15326_/D vssd1 vssd1 vccd1 vccd1 _15326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12538_ _12366_/A _12533_/X _12537_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12545_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15257_ _15258_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _12644_/A1 _12464_/X _12468_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12470_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14208_ _15364_/CLK _14208_/D vssd1 vssd1 vccd1 vccd1 _14208_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12797__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15188_ _15188_/CLK _15188_/D vssd1 vssd1 vccd1 vccd1 _15188_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07042__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ _15360_/CLK _14139_/D vssd1 vssd1 vccd1 vccd1 _14139_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout409 _07115_/Y vssd1 vssd1 vccd1 vccd1 _07131_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__12549__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _14036_/Q _06960_/Y _14026_/Q vssd1 vssd1 vccd1 vccd1 _06961_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08700_ _08776_/A _09860_/A _08573_/X _08574_/X _09858_/A vssd1 vssd1 vccd1 vccd1
+ _08705_/A sky130_fd_sc_hd__a32o_1
XANTENNA_hold2505_A _08250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _09679_/B _09824_/B _09679_/A vssd1 vssd1 vccd1 vccd1 _09681_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_158_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08631_ _08631_/A _12256_/A vssd1 vssd1 vccd1 vccd1 _08631_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08562_ hold777/A _14536_/Q _14696_/Q _14760_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08562_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_166_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12721__S0 _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ hold391/X _12329_/A _07528_/S vssd1 vssd1 vccd1 vccd1 hold392/A sky130_fd_sc_hd__mux2_1
XFILLER_0_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08493_ _08776_/B _08926_/A _08404_/X _08403_/X _09542_/A vssd1 vssd1 vccd1 vccd1
+ _08500_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15270_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07444_ _08253_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _14074_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12929__A1 _13398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07375_ _07364_/X _07374_/X _14051_/Q _12308_/A vssd1 vssd1 vccd1 vccd1 _07375_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09114_ _11320_/A _09114_/B vssd1 vssd1 vccd1 vccd1 _09114_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11887__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ _09045_/A _09167_/B _09045_/C vssd1 vssd1 vccd1 vccd1 _09047_/B sky130_fd_sc_hd__nand3_4
XANTENNA__10507__D _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13387__B _13387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 hold430/A vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12291__B _13468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 hold441/A vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10804__B _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 hold452/A vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold463 hold463/A vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10092__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold485 hold485/A vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold496/A vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13106__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09947_ _11497_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09947_/Y sky130_fd_sc_hd__nor2_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _10142_/A _10316_/B _09878_/C _10030_/A vssd1 vssd1 vccd1 vccd1 _10030_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _07776_/X vssd1 vssd1 vccd1 vccd1 _14392_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 _14461_/Q vssd1 vssd1 vccd1 vccd1 hold1141/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08533__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _08829_/A _08829_/B _08829_/C vssd1 vssd1 vccd1 vccd1 _08829_/Y sky130_fd_sc_hd__nor3_2
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 _11810_/X vssd1 vssd1 vccd1 vccd1 _14634_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 _15392_/Q vssd1 vssd1 vccd1 vccd1 hold1163/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 _11949_/X vssd1 vssd1 vccd1 vccd1 _14769_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 _14807_/Q vssd1 vssd1 vccd1 vccd1 hold1185/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1196 _11776_/X vssd1 vssd1 vccd1 vccd1 _14601_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ hold965/X _13727_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 hold966/A sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12617__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ hold1545/X _13691_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__mux2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _14958_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_178_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13510_ _13724_/A1 hold1937/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13510_/X sky130_fd_sc_hd__mux2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10719_/X _10720_/Y _10505_/Y _10548_/X vssd1 vssd1 vccd1 vccd1 _10722_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14490_ _15425_/CLK _14490_/D vssd1 vssd1 vccd1 vccd1 _14490_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _13459_/A _13441_/B vssd1 vssd1 vccd1 vccd1 _15214_/D sky130_fd_sc_hd__and2_1
X_10653_ _11594_/A _11588_/B _10457_/X _10456_/X _10283_/C vssd1 vssd1 vccd1 vccd1
+ _10658_/A sky130_fd_sc_hd__a32o_1
XANTENNA__13042__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _13373_/A _13372_/B vssd1 vssd1 vccd1 vccd1 _15163_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10584_ _11497_/A _10581_/X _10583_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _10585_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09261__A2 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ _15116_/CLK _15111_/D vssd1 vssd1 vccd1 vccd1 _15111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11797__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _12379_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and2_1
XFILLER_0_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07576__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ _15042_/CLK _15042_/D vssd1 vssd1 vccd1 vccd1 _15042_/Q sky130_fd_sc_hd__dfxtp_1
X_12254_ _12254_/A _12254_/B vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09644__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08447__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _11390_/A _11623_/A _11206_/C _11386_/A vssd1 vssd1 vccd1 vccd1 _11207_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08221__B1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12185_ hold2535/X _12195_/A2 _12184_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12185_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08772__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11136_ _11510_/A1 _11129_/Y _11131_/Y _11133_/Y _11135_/Y vssd1 vssd1 vccd1 vccd1
+ _11136_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_208_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13517__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _11067_/A _11240_/B _11067_/C vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__and3_2
XANTENNA__12856__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07515__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10129_/A _10827_/C _10019_/C _10019_/D vssd1 vssd1 vccd1 vccd1 _10020_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14826_ _14844_/CLK _14826_/D vssd1 vssd1 vccd1 vccd1 _14826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10882__A2 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11506__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14757_ _15398_/CLK _14757_/D vssd1 vssd1 vccd1 vccd1 _14757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12657__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11969_ hold1939/X _13724_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11969_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_137_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15062_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11561__A _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13708_ hold1469/X _13708_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13708_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14688_ _15397_/CLK hold720/X vssd1 vssd1 vccd1 vccd1 hold719/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13639_ _08179_/A _13625_/C _13638_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15352_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08292__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10608__C _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09788__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07160_ _13661_/A1 hold1523/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07160_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15309_ _15309_/CLK _15309_/D vssd1 vssd1 vccd1 vccd1 _15309_/Q sky130_fd_sc_hd__dfxtp_1
X_07091_ _13727_/A1 hold1729/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07091_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13336__A1 input153/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12544__C1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09801_ _15411_/Q _14546_/Q _14706_/Q _14770_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09801_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_157_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07993_ _08197_/A _07993_/B vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09732_ _09733_/A _09733_/B _09733_/C vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__o21a_2
X_06944_ _06944_/A vssd1 vssd1 vccd1 vccd1 _06944_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09663_ _09663_/A _09813_/B _09663_/C vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__and3_1
XFILLER_0_179_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08614_ _08614_/A _08614_/B vssd1 vssd1 vccd1 vccd1 _08616_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09594_ _09451_/X _09453_/Y _09592_/X _09593_/Y vssd1 vssd1 vccd1 vccd1 _09692_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08545_ _13558_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08545_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _14612_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout440_A _07512_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout538_A _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ _09816_/A _09712_/A vssd1 vssd1 vccd1 vccd1 _08476_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07160__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__B _12286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ _07427_/A _13317_/A vssd1 vssd1 vccd1 vccd1 _14057_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_135_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08126__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07358_ _07362_/D _07357_/X _07351_/A vssd1 vssd1 vccd1 vccd1 _07358_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08780__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13398__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14932__D _14932_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ _11623_/A _09724_/C vssd1 vssd1 vccd1 vccd1 _07290_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13327__A1 input149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _09027_/B _09027_/C _09027_/A vssd1 vssd1 vccd1 vccd1 _09030_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08203__B1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__B1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 _10304_/D vssd1 vssd1 vccd1 vccd1 _09864_/D sky130_fd_sc_hd__buf_4
XFILLER_0_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout751 _14951_/Q vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__buf_4
Xfanout762 _11561_/A vssd1 vssd1 vccd1 vccd1 _08809_/D sky130_fd_sc_hd__clkbuf_8
Xfanout773 _11333_/B vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__buf_4
X_13990_ _15296_/CLK _13990_/D vssd1 vssd1 vccd1 vccd1 _13990_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout784 _14942_/Q vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__buf_4
Xfanout795 _14491_/Q vssd1 vssd1 vccd1 vccd1 _12988_/C1 sky130_fd_sc_hd__buf_8
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12933__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ _14355_/Q hold567/A _12941_/S vssd1 vssd1 vccd1 vccd1 _12941_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10313__A1 _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12872_ hold793/A _14515_/Q _14643_/Q _14739_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12872_/X sky130_fd_sc_hd__mux4_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _15209_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _15035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ _15380_/CLK hold508/X vssd1 vssd1 vccd1 vccd1 hold507/A sky130_fd_sc_hd__dfxtp_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_133 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ hold1809/X hold2765/A _11828_/S vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15190_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_144 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_155 _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_177 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ _15439_/CLK hold694/X vssd1 vssd1 vccd1 vccd1 hold693/A sky130_fd_sc_hd__dfxtp_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10616__A2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_188 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ _13740_/A1 hold1487/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11754_/X sky130_fd_sc_hd__mux2_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_199 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07070__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10704_/B _10704_/C _10704_/A vssd1 vssd1 vccd1 vccd1 _10707_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07493__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14473_ _15276_/CLK hold874/X vssd1 vssd1 vccd1 vccd1 hold873/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ input45/X _13648_/B vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13424_ _13440_/S _13424_/B vssd1 vssd1 vccd1 vccd1 _13424_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10636_ _10819_/A _10635_/C _10635_/A vssd1 vssd1 vccd1 vccd1 _10673_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_181_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output192_A _15173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11041__A2 _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13355_ _13360_/A _13355_/B vssd1 vssd1 vccd1 vccd1 _15146_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12416__S _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ _11288_/A1 _10566_/Y _10435_/X vssd1 vssd1 vccd1 vccd1 _13456_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__13318__A1 input146/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _07437_/A _14031_/Q _14034_/Q _13240_/A vssd1 vssd1 vccd1 vccd1 _12306_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13101__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ input70/X fanout1/X _13285_/X vssd1 vssd1 vccd1 vccd1 _13287_/B sky130_fd_sc_hd__a21oi_1
X_10498_ _10498_/A _10498_/B _10498_/C vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__or3_4
X_15025_ _15188_/CLK _15025_/D vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12237_ _14622_/Q _14718_/Q _12237_/S vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__mux2_1
X_12168_ _14895_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__or2_1
XFILLER_0_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11119_ hold265/A hold531/A _14618_/Q _13987_/Q _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _11119_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12099_ hold2404/X _12099_/A2 _12098_/X _13499_/A vssd1 vssd1 vccd1 vccd1 _12099_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09026__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12924__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 dmemresp_rdata[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11990__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14809_ _15421_/CLK hold372/X vssd1 vssd1 vccd1 vccd1 hold371/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ _08329_/B _08329_/C _08329_/A vssd1 vssd1 vccd1 vccd1 _08331_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11804__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10619__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13006__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _13554_/B _08261_/B _08261_/C vssd1 vssd1 vccd1 vccd1 _08261_/X sky130_fd_sc_hd__or3_1
XFILLER_0_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13710__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__C _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ hold1451/X _13680_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 _07212_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08192_ _14788_/Q _14500_/Q _14628_/Q _14724_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08193_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08659__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _13744_/A1 hold2233/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07143_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13309__A1 input143/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10240__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _13679_/A1 hold1349/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput310 _14871_/Q vssd1 vssd1 vccd1 vccd1 out1[26] sky130_fd_sc_hd__buf_12
XFILLER_0_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput321 _14852_/Q vssd1 vssd1 vccd1 vccd1 out1[7] sky130_fd_sc_hd__buf_12
Xoutput332 _14830_/Q vssd1 vssd1 vccd1 vccd1 out2[17] sky130_fd_sc_hd__buf_12
XFILLER_0_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput343 _14840_/Q vssd1 vssd1 vccd1 vccd1 out2[27] sky130_fd_sc_hd__buf_12
XFILLER_0_168_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput354 _14821_/Q vssd1 vssd1 vccd1 vccd1 out2[8] sky130_fd_sc_hd__buf_12
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout390_A _11652_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _07976_/A _07976_/B vssd1 vssd1 vccd1 vccd1 _13345_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09581__D _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09715_ _09715_/A _09715_/B _09715_/C vssd1 vssd1 vccd1 vccd1 _09715_/Y sky130_fd_sc_hd__nand3_1
X_06927_ _14023_/Q vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__inv_2
XANTENNA_fanout655_A _15068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ _14673_/Q _13946_/Q hold915/A _13914_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09647_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_97_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06994__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09577_ _09575_/X _09577_/B vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14927__D _14927_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_A _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08528_ _08378_/A _08528_/B _09133_/A _08528_/D vssd1 vssd1 vccd1 vccd1 _08530_/D
+ sky130_fd_sc_hd__and4b_1
XANTENNA__08925__D _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08459_ hold965/A _13936_/Q hold765/A _13904_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08460_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_147_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11351__D _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ _11470_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _11471_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_6__f_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ _11504_/A _10418_/X _10420_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _10422_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12236__S _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ _13373_/A _13140_/B vssd1 vssd1 vccd1 vccd1 _15005_/D sky130_fd_sc_hd__nor2_1
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_131_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06986__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ hold953/A hold677/A hold451/A _14392_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _13071_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10283_ _11598_/A _11590_/A _10283_/C _11570_/B vssd1 vssd1 vccd1 vccd1 _10285_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12022_ _14984_/Q hold2656/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12022_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07935__C1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07065__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _10425_/S0 sky130_fd_sc_hd__buf_6
Xfanout581 _15218_/Q vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__clkbuf_8
Xfanout592 _09979_/D vssd1 vssd1 vccd1 vccd1 _11537_/B sky130_fd_sc_hd__clkbuf_8
X_13973_ _15371_/CLK _13973_/D vssd1 vssd1 vccd1 vccd1 _13973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09152__A1 _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__B1 _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ _13886_/Q _14014_/Q _13854_/Q _13822_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12924_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08685__A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _13080_/A1 _12854_/X _12852_/X vssd1 vssd1 vccd1 vccd1 _13161_/B sky130_fd_sc_hd__a21oi_4
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ hold569/X _13512_/A0 _11812_/S vssd1 vssd1 vccd1 vccd1 hold570/A sky130_fd_sc_hd__mux2_1
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12917_/A1 _12785_/X _12844_/A1 vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__a21o_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14557_/CLK hold440/X vssd1 vssd1 vccd1 vccd1 hold439/A sky130_fd_sc_hd__dfxtp_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _13657_/A1 hold2007/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13530__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14456_ _15390_/CLK _14456_/D vssd1 vssd1 vccd1 vccd1 _14456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11668_ _15052_/Q hold1157/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11668_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13407_ hold2354/X _13468_/A _13406_/Y _13409_/A vssd1 vssd1 vccd1 vccd1 _15197_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08851__C _08851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10619_ _11563_/A _11588_/B _10619_/C _10619_/D vssd1 vssd1 vccd1 vccd1 _10620_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14387_ _15383_/CLK _14387_/D vssd1 vssd1 vccd1 vccd1 _14387_/Q sky130_fd_sc_hd__dfxtp_1
X_11599_ _11599_/A _11599_/B vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10222__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13338_ _13338_/A _13338_/B vssd1 vssd1 vccd1 vccd1 _15132_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10773__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13269_ _13287_/A _13269_/B vssd1 vssd1 vccd1 vccd1 _15109_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _15268_/CLK _15008_/D vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13711__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10525__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2408 _14863_/Q vssd1 vssd1 vccd1 vccd1 hold2408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10525__B2 _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2419 _12095_/X vssd1 vssd1 vccd1 vccd1 _14859_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07830_ _12247_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07830_/Y sky130_fd_sc_hd__nor2_1
Xhold1707 _14252_/Q vssd1 vssd1 vccd1 vccd1 hold1707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1718 _07117_/X vssd1 vssd1 vccd1 vccd1 _13927_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10621__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1729 _13904_/Q vssd1 vssd1 vccd1 vccd1 hold1729/X sky130_fd_sc_hd__dlygate4sd3_1
X_07761_ _13666_/A1 hold1783/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07761_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_194_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09500_ hold217/A hold537/A hold613/A _13977_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09500_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13705__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10828__A2 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07692_ hold1285/X _13665_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 _07692_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08595__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08351__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _10142_/B _09430_/X _09429_/X vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2787_A _15102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09362_ _15376_/Q _15279_/Q hold689/A _14380_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09362_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_93_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09446__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08313_ _11340_/A _09437_/A _08312_/C _08312_/D vssd1 vssd1 vccd1 vccd1 _08314_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09293_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08244_ _08244_/A _08244_/B _08244_/C vssd1 vssd1 vccd1 vccd1 _08244_/X sky130_fd_sc_hd__and3_1
XFILLER_0_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_33 _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_44 _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_55 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_66 _15031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11005__A2 _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_77 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__S _12056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _13380_/B vssd1 vssd1 vccd1 vccd1 _08175_/Y sky130_fd_sc_hd__inv_2
XANTENNA_99 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12753__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07126_ _13727_/A1 hold2075/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07126_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10764__A1 _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ _13662_/A1 hold1823/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06989__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput162 _15165_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[0] sky130_fd_sc_hd__buf_12
XANTENNA__13702__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13395__B _13395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput173 _15166_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[1] sky130_fd_sc_hd__buf_12
Xoutput184 _15167_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[2] sky130_fd_sc_hd__buf_12
XANTENNA_fanout772_A _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 _06963_/X vssd1 vssd1 vccd1 vccd1 dmemreq_val sky130_fd_sc_hd__buf_12
XANTENNA__08489__B _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _07959_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07961_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_203_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09134__A1 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12364__S1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ _10970_/A _10970_/B _11150_/B vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07145__A0 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07613__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09629_ _15152_/Q _09925_/A2 _07390_/A vssd1 vssd1 vccd1 vccd1 _09629_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11643__B _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ hold969/A _14119_/Q _12641_/S vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_195_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11244__A2 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12571_ _15368_/Q _15271_/Q _15079_/Q _14372_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12571_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_109_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15422_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _14569_/CLK hold366/X vssd1 vssd1 vccd1 vccd1 hold365/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15290_ _15387_/CLK _15290_/D vssd1 vssd1 vccd1 vccd1 _15290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _15080_/CLK _14241_/D vssd1 vssd1 vccd1 vccd1 _14241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11453_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10275__A _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _10744_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__or2_1
XFILLER_0_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14172_ _15177_/CLK hold190/X vssd1 vssd1 vccd1 vccd1 _14172_/Q sky130_fd_sc_hd__dfxtp_1
X_11384_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10755__A1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ _13492_/A hold73/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__and2_1
X_10335_ _10336_/B _10336_/C _10336_/A vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _11287_/X _13104_/A2 _13053_/X vssd1 vssd1 vccd1 vccd1 _13054_/X sky130_fd_sc_hd__a21o_1
X_10266_ _10263_/C _10266_/B vssd1 vssd1 vccd1 vccd1 _10267_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ _12037_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _14815_/D sky130_fd_sc_hd__and2_1
XFILLER_0_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10197_ _10193_/Y _10194_/X _09987_/Y _09989_/X vssd1 vssd1 vccd1 vccd1 _10198_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_206_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13525__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13956_ _15068_/CLK _13956_/D vssd1 vssd1 vccd1 vccd1 _13956_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07523__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ _13171_/A _12907_/B vssd1 vssd1 vccd1 vccd1 _14964_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12680__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ _15382_/CLK _13887_/D vssd1 vssd1 vccd1 vccd1 _13887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09023__B _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12838_ _12917_/B1 hold2812/X _12837_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12845_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12769_ _12950_/S0 _12764_/X _12768_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12770_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15225_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14508_ _15184_/CLK hold670/X vssd1 vssd1 vccd1 vccd1 hold669/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 dmemresp_rdata[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10185__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput31 dmemresp_rdata[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
X_14439_ _15309_/CLK _14439_/D vssd1 vssd1 vccd1 vccd1 _14439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput42 imemresp_data[18] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 imemresp_data[28] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 imemresp_data[9] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
Xinput75 in0[19] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
Xhold804 hold804/A vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 in0[29] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_1
Xhold815 hold815/A vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold826 hold826/A vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 in1[0] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
Xhold837 hold837/A vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold848 hold848/A vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold2535_A _14999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13496__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ _10185_/A _11378_/C _09981_/C _10182_/A vssd1 vssd1 vccd1 vccd1 _09982_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold859 hold859/A vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08931_ _08930_/B _08930_/C _08930_/A vssd1 vssd1 vccd1 vccd1 _08932_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2205 _14226_/Q vssd1 vssd1 vccd1 vccd1 hold2205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2216 _11942_/X vssd1 vssd1 vccd1 vccd1 _14762_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08862_ _09087_/B _09087_/C vssd1 vssd1 vccd1 vccd1 _08862_/Y sky130_fd_sc_hd__xnor2_1
Xhold2227 _15070_/Q vssd1 vssd1 vccd1 vccd1 hold2227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2238 _11992_/X vssd1 vssd1 vccd1 vccd1 _14811_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1504 _07208_/X vssd1 vssd1 vccd1 vccd1 _14015_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2249 _13921_/Q vssd1 vssd1 vccd1 vccd1 hold2249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1515 _14628_/Q vssd1 vssd1 vccd1 vccd1 hold1515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _07153_/X vssd1 vssd1 vccd1 vccd1 _13961_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ hold275/A hold301/A _14591_/Q _13960_/Q _12198_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _07813_/X sky130_fd_sc_hd__mux4_1
X_08793_ _08908_/A _09026_/B _09712_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _08794_/C
+ sky130_fd_sc_hd__nand4_1
Xhold1537 _13808_/Q vssd1 vssd1 vccd1 vccd1 hold1537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1548 _07152_/X vssd1 vssd1 vccd1 vccd1 _13960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _14272_/Q vssd1 vssd1 vccd1 vccd1 hold1559/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07744_ _07744_/A _11729_/B _14090_/Q vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__or3_2
XANTENNA__12346__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11474__A2 _11474_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ hold1429/X _13714_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 _07675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ _09410_/X _09412_/Y _09305_/B _09307_/B vssd1 vssd1 vccd1 vccd1 _09414_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _09346_/B _09346_/C _09346_/A vssd1 vssd1 vccd1 vccd1 _09347_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout520_A _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout618_A _15205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15398_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _09275_/A _09275_/B _09146_/B vssd1 vssd1 vccd1 vccd1 _09277_/D sky130_fd_sc_hd__o21bai_1
XFILLER_0_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10807__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ _08226_/A _08226_/B _08226_/C vssd1 vssd1 vccd1 vccd1 _08228_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10526__C _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08158_ _08156_/B _08209_/B _08156_/A vssd1 vssd1 vccd1 vccd1 _08158_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ _13745_/A1 hold2135/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07109_/X sky130_fd_sc_hd__mux2_1
X_08089_ _08677_/A _11517_/A _08089_/C _08161_/B vssd1 vssd1 vccd1 vccd1 _08093_/A
+ sky130_fd_sc_hd__and4_2
XANTENNA__09961__A1_N _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10122_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07608__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15250_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09355__A1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _10050_/B _10050_/C _10050_/A vssd1 vssd1 vccd1 vccd1 _10052_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08012__B _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2750 _15173_/Q vssd1 vssd1 vccd1 vccd1 hold2750/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2761 _15107_/Q vssd1 vssd1 vccd1 vccd1 hold2761/X sky130_fd_sc_hd__buf_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2772 _15192_/Q vssd1 vssd1 vccd1 vccd1 hold2772/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2783 _15042_/Q vssd1 vssd1 vccd1 vccd1 hold2783/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2794 _15066_/Q vssd1 vssd1 vccd1 vccd1 hold2794/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _14569_/CLK _13810_/D vssd1 vssd1 vccd1 vccd1 _13810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12337__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _15270_/CLK hold666/X vssd1 vssd1 vccd1 vccd1 hold665/A sky130_fd_sc_hd__dfxtp_1
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__A2 _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09124__A _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ hold355/X _13741_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__mux2_1
X_10953_ _07299_/B _07302_/B _10077_/B _10952_/X _07297_/Y vssd1 vssd1 vccd1 vccd1
+ _10955_/A sky130_fd_sc_hd__a311o_1
XANTENNA__12662__A1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ hold447/X _13738_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold448/A sky130_fd_sc_hd__mux2_1
X_10884_ _10881_/X _10882_/Y _10639_/C _10641_/A vssd1 vssd1 vccd1 vccd1 _10885_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_195_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15411_ _15411_/CLK _15411_/D vssd1 vssd1 vccd1 vccd1 _15411_/Q sky130_fd_sc_hd__dfxtp_1
X_12623_ hold247/A hold365/A _14601_/Q _13970_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12623_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_156_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08682__B _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15427_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ _15422_/CLK _15342_/D vssd1 vssd1 vccd1 vccd1 _15342_/Q sky130_fd_sc_hd__dfxtp_2
X_12554_ _13383_/B _12325_/B _12553_/X vssd1 vssd1 vccd1 vccd1 _12554_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ hold367/A hold769/A hold535/A _14393_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11505_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07298__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15273_ _15440_/CLK _15273_/D vssd1 vssd1 vccd1 vccd1 _15273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12485_ _14660_/Q _13933_/Q _12491_/S vssd1 vssd1 vccd1 vccd1 _12485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09794__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14224_ _15449_/CLK _14224_/D vssd1 vssd1 vccd1 vccd1 _14224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _11146_/A _11146_/C _11146_/B vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11925__A0 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14155_ _15442_/CLK hold170/X vssd1 vssd1 vccd1 vccd1 _14155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11367_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07518__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13106_ _13106_/A1 _13171_/B _08637_/Y vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__o21a_1
X_10318_ _10318_/A _10483_/B _10318_/C vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__nand3_1
X_14086_ _15214_/CLK _14086_/D vssd1 vssd1 vccd1 vccd1 _14086_/Q sky130_fd_sc_hd__dfxtp_2
X_11298_ _11486_/B _11296_/Y _11297_/Y _13591_/A2 vssd1 vssd1 vccd1 vccd1 _11298_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13099_/S1 _13034_/X _13036_/X vssd1 vssd1 vccd1 vccd1 _13037_/X sky130_fd_sc_hd__a21o_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ hold425/A _14226_/Q hold467/A _14480_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10250_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08554__C1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09960__C _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11564__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_182_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14988_ _15248_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 _14988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12379__B _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _15440_/CLK _13939_/D vssd1 vssd1 vccd1 vccd1 _13939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07460_ _07460_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14090_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08873__A _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12405__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ _10233_/A _11650_/B vssd1 vssd1 vccd1 vccd1 _07391_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15325_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09130_ _09714_/A _10126_/A _10126_/B _09571_/A vssd1 vssd1 vccd1 vccd1 _09130_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10416__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__A2 _13165_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_77_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _09060_/A _09060_/B _09021_/Y vssd1 vssd1 vccd1 vccd1 _09061_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_120_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ _08312_/A _08012_/B _08012_/C _08012_/D vssd1 vssd1 vccd1 vccd1 _08014_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold601 hold601/A vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 hold612/A vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08388__A2 _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold623 hold623/A vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold634 hold634/A vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10643__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 hold645/A vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 hold656/A vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 hold667/A vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09963_ _09963_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__or2_1
XANTENNA__09209__A _13390_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold678 hold678/A vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 hold689/A vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_135_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08914_ _08914_/A _08914_/B vssd1 vssd1 vccd1 vccd1 _08915_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2002 _07169_/X vssd1 vssd1 vccd1 vccd1 _13977_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2013 _14367_/Q vssd1 vssd1 vccd1 vccd1 hold2013/X sky130_fd_sc_hd__dlygate4sd3_1
X_09894_ _10052_/A _09894_/B _09741_/A vssd1 vssd1 vccd1 vccd1 _09896_/C sky130_fd_sc_hd__nor3b_4
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 _11704_/X vssd1 vssd1 vccd1 vccd1 _14500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2035 _14775_/Q vssd1 vssd1 vccd1 vccd1 hold2035/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 _13846_/Q vssd1 vssd1 vccd1 vccd1 hold1301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2046 _07043_/X vssd1 vssd1 vccd1 vccd1 _13860_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08846_/B _08846_/C _07323_/B vssd1 vssd1 vccd1 vccd1 _08845_/X sky130_fd_sc_hd__a21bo_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 _13901_/Q vssd1 vssd1 vccd1 vccd1 hold2057/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1312 _07670_/X vssd1 vssd1 vccd1 vccd1 _14291_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 _15398_/Q vssd1 vssd1 vccd1 vccd1 hold1323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12892__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2068 _11698_/X vssd1 vssd1 vccd1 vccd1 _14494_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout470_A _12128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2079 _13974_/Q vssd1 vssd1 vccd1 vccd1 hold2079/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _13687_/X vssd1 vssd1 vccd1 vccd1 _15393_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1345 _14391_/Q vssd1 vssd1 vccd1 vccd1 hold1345/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout568_A _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07994__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1356 _13504_/X vssd1 vssd1 vccd1 vccd1 _15262_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12319__S1 _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _08776_/A _08776_/B _09858_/B vssd1 vssd1 vccd1 vccd1 _08776_/X sky130_fd_sc_hd__and3_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1367 _14241_/Q vssd1 vssd1 vccd1 vccd1 hold1367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1378 _11974_/X vssd1 vssd1 vccd1 vccd1 _14793_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07163__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12289__B _13464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1389 _14780_/Q vssd1 vssd1 vccd1 vccd1 hold1389/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ hold539/X _13700_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold540/A sky130_fd_sc_hd__mux2_1
XANTENNA__12644__A1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__B1 _08773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10655__B1 _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ hold1273/X _13730_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 _07658_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14935__D _14935_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07589_ _13728_/A1 hold1665/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07589_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12509__S _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09328_ _09328_/A _09328_/B _09328_/C vssd1 vssd1 vccd1 vccd1 _09328_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_118_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08076__A1 _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08076__B2 _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _09257_/X _09259_/B vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_106_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07823__A1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09025__B1 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12270_ _13150_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _14919_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _11220_/A _11220_/B _11331_/B _11220_/D vssd1 vssd1 vccd1 vccd1 _11221_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__10186__A2 _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _11598_/A _11573_/B _14966_/Q _11597_/A vssd1 vssd1 vccd1 vccd1 _11155_/C
+ sky130_fd_sc_hd__a22o_1
X_10103_ _11510_/A1 _10096_/Y _10098_/Y _10100_/Y _10102_/Y vssd1 vssd1 vccd1 vccd1
+ _10103_/X sky130_fd_sc_hd__o32a_1
XANTENNA__12558__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ _11082_/A _11082_/B _11082_/C vssd1 vssd1 vccd1 vccd1 _11086_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11135__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _10142_/B _10316_/B _10035_/C _10141_/A vssd1 vssd1 vccd1 vccd1 _10036_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08000__A1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ _15416_/CLK _14911_/D vssd1 vssd1 vccd1 vccd1 _14911_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__B _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2580 _15135_/Q vssd1 vssd1 vccd1 vccd1 hold2580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _14842_/CLK _14842_/D vssd1 vssd1 vccd1 vccd1 _14842_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2591 _14993_/Q vssd1 vssd1 vccd1 vccd1 hold2591/X sky130_fd_sc_hd__buf_2
XFILLER_0_76_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07073__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1890 _07053_/X vssd1 vssd1 vccd1 vccd1 _13869_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ hold1231/X _13674_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__mux2_1
X_14773_ _15408_/CLK _14773_/D vssd1 vssd1 vccd1 vccd1 _14773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13724_ hold1655/X _13724_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 _13724_/X sky130_fd_sc_hd__mux2_1
X_10936_ _11504_/A _10933_/X _10935_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _10937_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07801__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ _10866_/A _10866_/B _10866_/C vssd1 vssd1 vccd1 vccd1 _10868_/B sky130_fd_sc_hd__a21oi_1
X_13655_ hold949/X _13655_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold950/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09301__B _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12606_ _13081_/A1 _13151_/B _08637_/Y vssd1 vssd1 vccd1 vccd1 _12607_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08067__A1 _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A _13586_/B vssd1 vssd1 vccd1 vccd1 _13586_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _11594_/A _11563_/A _11606_/B _11570_/B vssd1 vssd1 vccd1 vccd1 _10801_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__10949__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10447__B _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15325_ _15325_/CLK _15325_/D vssd1 vssd1 vccd1 vccd1 _15325_/Q sky130_fd_sc_hd__dfxtp_1
X_12537_ _12668_/A1 _12534_/X _12536_/X vssd1 vssd1 vccd1 vccd1 _12537_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__C _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12468_ _12343_/A _12465_/X _12467_/X vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12246__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15256_ _15256_/CLK hold110/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09567__A1 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ _11551_/A _11418_/C _11418_/A vssd1 vssd1 vccd1 vccd1 _11420_/C sky130_fd_sc_hd__a21o_1
X_14207_ _14754_/CLK _14207_/D vssd1 vssd1 vccd1 vccd1 _14207_/Q sky130_fd_sc_hd__dfxtp_1
X_15187_ _15278_/CLK _15187_/D vssd1 vssd1 vccd1 vccd1 _15187_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12797__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ _13865_/Q hold681/A _13833_/Q _13801_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12399_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ _15390_/CLK hold392/X vssd1 vssd1 vccd1 vccd1 hold391/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11993__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ _14028_/Q _14036_/Q vssd1 vssd1 vccd1 vccd1 _06960_/Y sky130_fd_sc_hd__nor2_1
X_14069_ _15222_/CLK _14069_/D vssd1 vssd1 vccd1 vccd1 _14069_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12549__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15364_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11126__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08630_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _08630_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ _08989_/A _08561_/B vssd1 vssd1 vccd1 vccd1 _08561_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13713__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07512_ _13716_/A _07644_/A vssd1 vssd1 vccd1 vccd1 _07512_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_18_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08492_ _08492_/A _08492_/B vssd1 vssd1 vccd1 vccd1 _08507_/A sky130_fd_sc_hd__and2_1
XANTENNA__12721__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07711__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07443_ _08179_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _14073_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__A1 _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12929__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07374_ _07370_/X _07371_/Y _07372_/X _07373_/Y _07369_/X vssd1 vssd1 vccd1 vccd1
+ _07374_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09113_ _09098_/Y _09103_/Y _09112_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09114_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09044_ _10185_/A _10022_/B _09043_/C _09167_/A vssd1 vssd1 vccd1 vccd1 _09045_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07947__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold420 hold420/A vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold431 hold431/A vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold442 hold442/A vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10804__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold453 hold453/A vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold464 hold464/A vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold475/A vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold486 hold486/A vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold497 hold497/A vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06997__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ hold593/A _14224_/Q hold691/A hold729/A _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _09947_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11117__A1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _10142_/A _10316_/B _09878_/C _10030_/A vssd1 vssd1 vccd1 vccd1 _09879_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout852_A _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _13738_/X vssd1 vssd1 vccd1 vccd1 _15448_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 _14306_/Q vssd1 vssd1 vccd1 vccd1 hold1131/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _11658_/X vssd1 vssd1 vccd1 vccd1 _14461_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _08824_/X _08826_/Y _08717_/B _08717_/Y vssd1 vssd1 vccd1 vccd1 _08829_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 _13994_/Q vssd1 vssd1 vccd1 vccd1 hold1153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 _13686_/X vssd1 vssd1 vccd1 vccd1 _15392_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1175 _15360_/Q vssd1 vssd1 vccd1 vccd1 hold1175/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _11988_/X vssd1 vssd1 vccd1 vccd1 _14807_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _08989_/A _08756_/X _08758_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08760_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12617__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1197 _14914_/Q vssd1 vssd1 vccd1 vccd1 _13475_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11770_ hold1949/X _13657_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11770_/X sky130_fd_sc_hd__mux2_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07621__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10721_ _10505_/Y _10548_/X _10719_/X _10720_/Y vssd1 vssd1 vccd1 vccd1 _10721_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _09346_/A _12277_/B _13440_/S vssd1 vssd1 vccd1 vccd1 _13441_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13042__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13371_ _13373_/A _13371_/B vssd1 vssd1 vccd1 vccd1 _15162_/D sky130_fd_sc_hd__nor2_1
X_10583_ _11507_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__or2_1
XFILLER_0_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15110_ _15116_/CLK _15110_/D vssd1 vssd1 vccd1 vccd1 _15110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12322_ _12601_/A _12321_/X _12294_/X vssd1 vssd1 vccd1 vccd1 _12322_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__13578__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12228__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15041_ _15434_/CLK _15041_/D vssd1 vssd1 vccd1 vccd1 _15041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12253_ hold2646/X input12/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13173_/B sky130_fd_sc_hd__mux2_2
XANTENNA__10283__A _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__B _07576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11204_ _11409_/A _11588_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11386_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__09644__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07068__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__A1 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ _14903_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__or2_1
XANTENNA__08221__B2 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11135_ _11493_/A _11134_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _11135_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07980__B1 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11066_ _11240_/A _11065_/C _11065_/A vssd1 vssd1 vccd1 vccd1 _11067_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12400__S0 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _10126_/A _10126_/B _11168_/A _11606_/A vssd1 vssd1 vccd1 vccd1 _10019_/D
+ sky130_fd_sc_hd__nand4_4
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12003__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14842_/CLK _14825_/D vssd1 vssd1 vccd1 vccd1 _14825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13533__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__A1 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _15361_/CLK _14756_/D vssd1 vssd1 vccd1 vccd1 _14756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11968_ hold1053/X _13657_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11968_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07531__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11561__B _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ hold679/X _13740_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold680/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10919_ _11288_/A1 _10918_/X _10778_/X vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__a21oi_4
X_14687_ _15429_/CLK _14687_/D vssd1 vssd1 vccd1 vccd1 _14687_/Q sky130_fd_sc_hd__dfxtp_1
X_11899_ _13654_/A1 hold2219/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13638_ input51/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__or2_1
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09788__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11988__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10608__D _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ _09213_/B _08441_/B _13568_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13569_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12792__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15308_ _15309_/CLK _15308_/D vssd1 vssd1 vccd1 vccd1 _15308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ _13693_/A1 hold2063/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11289__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15239_ _15244_/CLK hold124/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08748__C1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09800_ _10426_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09800_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13708__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07992_ hold603/A _14238_/Q hold779/A _14110_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _07993_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07706__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _09731_/A _09731_/B vssd1 vssd1 vccd1 vccd1 _09733_/C sky130_fd_sc_hd__xnor2_1
X_06943_ _06943_/A vssd1 vssd1 vccd1 vccd1 _06943_/Y sky130_fd_sc_hd__inv_6
XFILLER_0_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09662_ _09527_/A _09527_/B _09527_/C vssd1 vssd1 vccd1 vccd1 _09663_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08613_ _08614_/A _08614_/B vssd1 vssd1 vccd1 vccd1 _08613_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09593_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _13558_/A _14434_/Q _08544_/C vssd1 vssd1 vccd1 vccd1 _08856_/C sky130_fd_sc_hd__and3_1
XANTENNA__11283__A0 hold2779/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _09816_/A _08685_/C _08395_/D _08392_/X vssd1 vssd1 vccd1 vccd1 _08487_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout433_A _07778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07426_ _07426_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14056_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12458__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ _15340_/Q _15339_/Q _15331_/Q _15330_/Q vssd1 vssd1 vccd1 vccd1 _07357_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09876__B _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13398__B _13398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ _10827_/D _09724_/C vssd1 vssd1 vccd1 vccd1 _09205_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09027_ _09027_/A _09027_/B _09027_/C vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08203__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 _14958_/Q vssd1 vssd1 vccd1 vccd1 _11588_/B sky130_fd_sc_hd__clkbuf_8
Xfanout741 _10304_/D vssd1 vssd1 vccd1 vccd1 _09714_/D sky130_fd_sc_hd__buf_2
XANTENNA__07616__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout752 _11614_/A vssd1 vssd1 vccd1 vccd1 _10126_/B sky130_fd_sc_hd__buf_4
XANTENNA__12838__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _09778_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__nand2b_1
Xfanout763 _14948_/Q vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__clkbuf_8
Xfanout774 _11333_/B vssd1 vssd1 vccd1 vccd1 _09026_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout785 _14942_/Q vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__clkbuf_8
Xfanout796 _12366_/A vssd1 vssd1 vccd1 vccd1 _12642_/B1 sky130_fd_sc_hd__buf_6
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08062__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12940_ hold547/A _14131_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12940_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10313__A2 _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12871_ hold551/A hold951/A hold837/A _14384_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12871_/X sky130_fd_sc_hd__mux4_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _12284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _15379_/CLK _14610_/D vssd1 vssd1 vccd1 vccd1 _14610_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ hold295/X _11921_/A0 _11828_/S vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__mux2_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_145 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_167 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_178 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ _15056_/CLK _14541_/D vssd1 vssd1 vccd1 vccd1 _14541_/Q sky130_fd_sc_hd__dfxtp_1
X_11753_ _13739_/A1 hold1877/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__mux2_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10278__A _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_189 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/A _10704_/B _10704_/C vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__nand3_2
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11684_ _13715_/A1 hold1271/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11684_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14472_ _14472_/CLK _14472_/D vssd1 vssd1 vccd1 vccd1 _14472_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12449__S0 _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10635_ _10635_/A _10819_/A _10635_/C vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_126_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13423_ _08345_/B _13450_/A _13422_/Y _13178_/A vssd1 vssd1 vccd1 vccd1 _15205_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13354_ _13360_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _15145_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ _10436_/Y _10437_/X _10565_/X vssd1 vssd1 vccd1 vccd1 _10566_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output185_A _15195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12305_ _12294_/A _14035_/Q _12303_/X _12304_/X _15293_/Q vssd1 vssd1 vccd1 vccd1
+ _12308_/C sky130_fd_sc_hd__o2111a_1
XFILLER_0_84_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13285_ input134/X fanout6/X fanout4/X input102/X vssd1 vssd1 vccd1 vccd1 _13285_/X
+ sky130_fd_sc_hd__a22o_1
X_10497_ _10496_/A _10496_/B _10482_/Y vssd1 vssd1 vccd1 vccd1 _10498_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_121_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15024_ _15188_/CLK _15024_/D vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__dfxtp_1
X_12236_ _14782_/Q _14494_/Q _12237_/S vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12621__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09942__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12167_ hold2439/X _12173_/A2 _12166_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12167_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07526__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ _11113_/A _13591_/A2 _11104_/X _11117_/Y _13459_/A vssd1 vssd1 vccd1 vccd1
+ _11118_/X sky130_fd_sc_hd__o221a_1
X_12098_ _14989_/Q _12128_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12098_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12829__A1 _13394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09026__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ _11049_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12924__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 dmemresp_rdata[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14808_ _14926_/CLK hold564/X vssd1 vssd1 vccd1 vccd1 hold563/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09042__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08356__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14739_ _15372_/CLK _14739_/D vssd1 vssd1 vccd1 vccd1 _14739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08260_ _09494_/A1 _08258_/Y _08259_/X _09925_/A2 _15140_/Q vssd1 vssd1 vccd1 vccd1
+ _08261_/C sky130_fd_sc_hd__a32o_1
XFILLER_0_184_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13006__A1 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07211_ hold293/X _13679_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__mux2_1
XANTENNA__10338__D _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13499__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ hold647/A _15268_/Q _15076_/Q _14369_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08191_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07142_ _13743_/A1 hold1571/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07142_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10240__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07073_ _13744_/A1 hold1337/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput300 _14862_/Q vssd1 vssd1 vccd1 vccd1 out1[17] sky130_fd_sc_hd__buf_12
XFILLER_0_70_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput311 _14872_/Q vssd1 vssd1 vccd1 vccd1 out1[27] sky130_fd_sc_hd__buf_12
XFILLER_0_113_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12517__B1 _14490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput322 _14853_/Q vssd1 vssd1 vccd1 vccd1 out1[8] sky130_fd_sc_hd__buf_12
Xoutput333 _14831_/Q vssd1 vssd1 vccd1 vccd1 out2[18] sky130_fd_sc_hd__buf_12
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput344 _14841_/Q vssd1 vssd1 vccd1 vccd1 out2[28] sky130_fd_sc_hd__buf_12
XFILLER_0_140_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput355 _14822_/Q vssd1 vssd1 vccd1 vccd1 out2[9] sky130_fd_sc_hd__buf_12
XFILLER_0_168_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12342__S _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07944__B1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07975_ _07975_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _07976_/B sky130_fd_sc_hd__and2_1
XANTENNA__08121__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout383_A _11895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09714_ _09714_/A _09864_/A _09714_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09715_/C
+ sky130_fd_sc_hd__nand4_1
X_06926_ _06926_/A vssd1 vssd1 vccd1 vccd1 _06926_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07960__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _10426_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout550_A _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout648_A _15198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09576_ _09573_/Y _09574_/X _09434_/X _09436_/X vssd1 vssd1 vccd1 vccd1 _09577_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07171__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _09133_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08530_/C sky130_fd_sc_hd__nor2_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10098__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout815_A _14489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09887__A _09888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _12247_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08458_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08791__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07409_ _13501_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _14039_/D sky130_fd_sc_hd__and2_1
XFILLER_0_80_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08389_ _08389_/A _08389_/B _08389_/C vssd1 vssd1 vccd1 vccd1 _08393_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11559__A1 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10826__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _11493_/A _10420_/B vssd1 vssd1 vccd1 vccd1 _10420_/X sky130_fd_sc_hd__or2_1
XANTENNA__13202__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12756__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _10351_/A _15221_/Q vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13070_ _13070_/A _13070_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__or3b_1
X_10282_ _10282_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__xor2_2
X_12021_ _12059_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _14823_/D sky130_fd_sc_hd__and2_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10090__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _08763_/S0 vssd1 vssd1 vccd1 vccd1 _08868_/S0 sky130_fd_sc_hd__buf_8
Xfanout571 _11316_/S0 vssd1 vssd1 vccd1 vccd1 _11306_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_205_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout582 _15218_/Q vssd1 vssd1 vccd1 vccd1 _10338_/D sky130_fd_sc_hd__buf_2
Xfanout593 _09979_/D vssd1 vssd1 vccd1 vccd1 _10830_/B sky130_fd_sc_hd__clkbuf_4
X_13972_ _15367_/CLK _13972_/D vssd1 vssd1 vccd1 vccd1 _13972_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09152__A2 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ hold279/X hold297/A hold311/A _13982_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12923_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_38_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08685__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12854_ _13395_/B _13104_/A2 _12853_/X vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__a21o_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07081__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ hold375/X _13659_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold376/A sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12444__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ hold721/A _13945_/Q _12791_/S vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__mux2_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08112__B1 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11798__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _15389_/CLK hold386/X vssd1 vssd1 vccd1 vccd1 hold385/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ _13689_/A1 hold2239/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__mux2_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10470__A1 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14455_ _15325_/CLK _14455_/D vssd1 vssd1 vccd1 vccd1 _14455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11667_ _13698_/A1 hold1555/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ _13468_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13406_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10618_ _11563_/A _11588_/B _10619_/C _10619_/D vssd1 vssd1 vccd1 vccd1 _10620_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11598_ _11598_/A _14967_/Q vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08206__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14386_ _15093_/CLK _14386_/D vssd1 vssd1 vccd1 vccd1 _14386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13337_ input89/X fanout2/X _13336_/X vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__a21oi_1
X_10549_ _10548_/A _10548_/B _10548_/C _10548_/D vssd1 vssd1 vccd1 vccd1 _10549_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12951__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ input95/X fanout1/X _13267_/X vssd1 vssd1 vccd1 vccd1 _13269_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11567__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ _15177_/CLK _15007_/D vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09376__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12219_ _12252_/A _12252_/B _12219_/C _12219_/D vssd1 vssd1 vccd1 vccd1 _12219_/X
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__10471__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13199_ _13404_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _15064_/D sky130_fd_sc_hd__and2_1
Xhold2409 _12103_/X vssd1 vssd1 vccd1 vccd1 _14863_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10525__A2 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1708 _07629_/X vssd1 vssd1 vccd1 vccd1 _14252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 _15410_/Q vssd1 vssd1 vccd1 vccd1 hold1719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10621__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _13665_/A1 hold1371/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07760_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07691_ hold1499/X _13664_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 _07691_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08595__B _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ _10022_/A _11586_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _09430_/X sky130_fd_sc_hd__and3_1
XFILLER_0_189_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ _10244_/A _09358_/X _09360_/X vssd1 vssd1 vccd1 vccd1 _09361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08103__B1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ _08312_/A _09437_/A _08312_/C _08312_/D vssd1 vssd1 vccd1 vccd1 _08314_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13721__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12986__B1 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09292_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08243_ _08242_/B _08243_/B vssd1 vssd1 vccd1 vccd1 _08243_/X sky130_fd_sc_hd__and2b_1
XANTENNA_23 _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _14928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_45 _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_67 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08174_ _08173_/X _08174_/B vssd1 vssd1 vccd1 vccd1 _13380_/B sky130_fd_sc_hd__and2b_4
XFILLER_0_16_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_78 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_89 _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07125_ _13693_/A1 hold1979/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07056_ _13661_/A1 hold1421/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07056_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout598_A _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 _15175_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[10] sky130_fd_sc_hd__buf_12
Xoutput174 _15185_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[20] sky130_fd_sc_hd__buf_12
XFILLER_0_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput185 _15195_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[30] sky130_fd_sc_hd__buf_12
XANTENNA__07166__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput196 _14170_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[0] sky130_fd_sc_hd__buf_12
XFILLER_0_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11196__B _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07958_ _07958_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_199_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06909_ _15344_/Q vssd1 vssd1 vccd1 vccd1 _06909_/Y sky130_fd_sc_hd__inv_2
X_07889_ _08677_/A _11566_/A _07889_/C vssd1 vssd1 vccd1 vccd1 _07958_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09628_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _13361_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09559_ _09417_/B _09418_/Y _09557_/X _09558_/Y vssd1 vssd1 vccd1 vccd1 _09602_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_66_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12620__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _12570_/A _12570_/B _12601_/A vssd1 vssd1 vccd1 vccd1 _12577_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11452_ _11607_/B _11450_/X _11183_/A _11183_/Y vssd1 vssd1 vccd1 vccd1 _11453_/B
+ sky130_fd_sc_hd__a211o_1
X_14240_ _15428_/CLK hold914/X vssd1 vssd1 vccd1 vccd1 hold913/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08026__A _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__B _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ _09930_/A _10401_/X _10402_/X vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__o21ba_1
X_14171_ _15177_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _14171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12770__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11383_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10755__A2 _12286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _10333_/B _10333_/C _10333_/A vssd1 vssd1 vccd1 vccd1 _10336_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_131_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13122_ _13491_/A hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__and2_1
XFILLER_0_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _13746_/A1 _13103_/A2 _13078_/B1 _13201_/B vssd1 vssd1 vccd1 vccd1 _13053_/X
+ sky130_fd_sc_hd__a22o_1
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12004_ hold2548/X hold2708/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07076__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _10198_/B vssd1 vssd1 vccd1 vccd1 _10196_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_121_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12710__S _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08696__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout390 _11652_/Y vssd1 vssd1 vccd1 vccd1 _11684_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07804__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13955_ _15456_/CLK _13955_/D vssd1 vssd1 vccd1 vccd1 _13955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12906_ _13106_/A1 _13163_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12011__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13886_ _15093_/CLK _13886_/D vssd1 vssd1 vccd1 vccd1 _13886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08884__B2 _13186_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12939_/S1 _12834_/X _12836_/X vssd1 vssd1 vccd1 vccd1 _12837_/X sky130_fd_sc_hd__a21o_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12768_ _06942_/A _12765_/X _12767_/X vssd1 vssd1 vccd1 vccd1 _12768_/X sky130_fd_sc_hd__a21o_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__A _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14731_/CLK _14507_/D vssd1 vssd1 vccd1 vccd1 _14507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11640__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ hold1225/X _13673_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12699_ _13877_/Q hold713/A _13845_/Q _13813_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12699_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 dmemresp_rdata[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
X_14438_ _15309_/CLK _14438_/D vssd1 vssd1 vccd1 vccd1 _14438_/Q sky130_fd_sc_hd__dfxtp_1
Xinput21 dmemresp_rdata[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10185__B _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput32 dmemresp_rdata[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 imemresp_data[19] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput54 imemresp_data[29] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput65 in0[0] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold805 hold805/A vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _15365_/CLK _14369_/D vssd1 vssd1 vccd1 vccd1 _14369_/Q sky130_fd_sc_hd__dfxtp_1
Xinput76 in0[1] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold816 hold816/A vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 in0[2] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_1
Xinput98 in1[10] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
Xhold827 hold827/A vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold838 hold838/A vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 hold849/A vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _08930_/A _08930_/B _08930_/C vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2206 _07602_/X vssd1 vssd1 vccd1 vccd1 _14226_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2217 _13799_/Q vssd1 vssd1 vccd1 vccd1 hold2217/X sky130_fd_sc_hd__dlygate4sd3_1
X_08861_ _08856_/A _09222_/B _08860_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _08861_/X
+ sky130_fd_sc_hd__o211a_1
Xhold2228 _13206_/X vssd1 vssd1 vccd1 vccd1 _15070_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2239 _14530_/Q vssd1 vssd1 vccd1 vccd1 hold2239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1505 _14610_/Q vssd1 vssd1 vccd1 vccd1 hold1505/X sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07812_/X sky130_fd_sc_hd__or2_1
Xhold1516 _11804_/X vssd1 vssd1 vccd1 vccd1 _14628_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08792_ _09026_/B _09712_/A _09708_/B _08908_/A vssd1 vssd1 vccd1 vccd1 _08794_/B
+ sky130_fd_sc_hd__a22o_1
Xhold1527 _14118_/Q vssd1 vssd1 vccd1 vccd1 hold1527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 _06989_/X vssd1 vssd1 vccd1 vccd1 _13808_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 _13910_/Q vssd1 vssd1 vccd1 vccd1 hold1549/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09116__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _14088_/Q _14089_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _13502_/B sky130_fd_sc_hd__and3_2
XFILLER_0_197_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ hold813/X _15066_/Q _07676_/S vssd1 vssd1 vccd1 vccd1 hold814/A sky130_fd_sc_hd__mux2_1
XFILLER_0_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09413_ _09305_/B _09307_/B _09410_/X _09412_/Y vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11306__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ _09344_/A _09344_/B vssd1 vssd1 vccd1 vccd1 _09346_/C sky130_fd_sc_hd__and2_1
XFILLER_0_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09230__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09275_ _09275_/A _09275_/B _09146_/B vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout513_A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08226_ _08226_/A _08226_/B _08226_/C vssd1 vssd1 vccd1 vccd1 _08228_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12187__A1 _12120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08156_/B _08209_/B _08156_/A vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10526__D _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07108_ _13744_/A1 hold2249/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07108_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08088_ _10873_/A _09138_/A _08161_/A _08088_/D vssd1 vssd1 vccd1 vccd1 _08161_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_28_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout882_A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07039_ hold1657/X hold2765/A _07044_/S vssd1 vssd1 vccd1 vccd1 _07039_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13687__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10050_ _10050_/A _10050_/B _10050_/C vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09355__A2 _12277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__B1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2740 _14967_/Q vssd1 vssd1 vccd1 vccd1 _07295_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2751 _15128_/Q vssd1 vssd1 vccd1 vccd1 hold2751/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2762 _15116_/Q vssd1 vssd1 vccd1 vccd1 hold2762/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2773 _15121_/Q vssd1 vssd1 vccd1 vccd1 hold2773/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07624__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2784 _15132_/Q vssd1 vssd1 vccd1 vccd1 hold2784/X sky130_fd_sc_hd__buf_1
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2795 _15119_/Q vssd1 vssd1 vccd1 vccd1 hold2795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ hold329/X _13740_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__mux2_1
XFILLER_0_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10952_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10952_/X sky130_fd_sc_hd__or2_1
XANTENNA__11373__C _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13671_ hold377/X _13671_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold378/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10883_ _10639_/C _10641_/A _10881_/X _10882_/Y vssd1 vssd1 vccd1 vccd1 _10885_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_35_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15410_ _15410_/CLK _15410_/D vssd1 vssd1 vccd1 vccd1 _15410_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _14793_/Q _14505_/Q _14633_/Q _14729_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12622_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_195_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15341_ _15422_/CLK _15341_/D vssd1 vssd1 vccd1 vccd1 _15341_/Q sky130_fd_sc_hd__dfxtp_2
X_12553_ _13512_/A0 _12329_/B _12953_/B1 _13181_/B vssd1 vssd1 vccd1 vccd1 _12553_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10286__A _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _11504_/A _11504_/B vssd1 vssd1 vccd1 vccd1 _11504_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15272_ _15369_/CLK hold706/X vssd1 vssd1 vccd1 vccd1 hold705/A sky130_fd_sc_hd__dfxtp_1
X_12484_ _15434_/Q _13901_/Q _12491_/S vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14223_ _15448_/CLK _14223_/D vssd1 vssd1 vccd1 vccd1 _14223_/Q sky130_fd_sc_hd__dfxtp_1
X_11435_ _11435_/A _11435_/B vssd1 vssd1 vccd1 vccd1 _11443_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11366_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11366_/X sky130_fd_sc_hd__and2_1
XFILLER_0_105_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14154_ _14472_/CLK _14154_/D vssd1 vssd1 vccd1 vccd1 _14154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10317_ _11569_/A _10316_/B _10483_/A _10316_/D vssd1 vssd1 vccd1 vccd1 _10318_/C
+ sky130_fd_sc_hd__a22o_1
X_13105_ _12327_/A _13104_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _13171_/B sky130_fd_sc_hd__a21oi_1
X_14085_ _14105_/CLK _14085_/D vssd1 vssd1 vccd1 vccd1 _14085_/Q sky130_fd_sc_hd__dfxtp_1
X_11297_ _11297_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11297_/Y sky130_fd_sc_hd__nand2_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10248_ _15424_/Q _10248_/B vssd1 vssd1 vccd1 vccd1 _10248_/Y sky130_fd_sc_hd__nor2_1
X_13036_ _13092_/A1 _13035_/X _13100_/S0 vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_206_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12350__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _14941_/Q _15220_/Q _10180_/A vssd1 vssd1 vccd1 vccd1 _10179_/X sky130_fd_sc_hd__and3_1
XANTENNA__12440__S _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09960__D _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07534__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11564__B _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12638__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14987_ _14987_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _14987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12379__C _13376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13938_ _15372_/CLK _13938_/D vssd1 vssd1 vccd1 vccd1 _13938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12653__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13869_ _15040_/CLK _13869_/D vssd1 vssd1 vccd1 vccd1 _13869_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12676__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ _07390_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _07926_/A sky130_fd_sc_hd__nor2_2
XANTENNA__13063__C1 _14491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10416__A1 _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _09060_/A _09060_/B _09021_/Y vssd1 vssd1 vccd1 vccd1 _09060_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_0_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12169__A1 _12102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08011_ _08010_/B _08010_/C _08010_/A vssd1 vssd1 vccd1 vccd1 _08012_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_60_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12615__S _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10924__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold602 hold602/A vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07709__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 hold613/A vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 hold624/A vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold635 hold635/A vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10643__B _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 hold646/A vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold657 hold657/A vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 hold668/A vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _09959_/Y _10170_/A _11335_/A _10338_/C vssd1 vssd1 vccd1 vccd1 _10170_/B
+ sky130_fd_sc_hd__and4bb_1
Xhold679 hold679/A vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08913_ _08912_/A _08912_/B _08912_/C vssd1 vssd1 vccd1 vccd1 _08914_/B sky130_fd_sc_hd__a21oi_1
Xhold2003 _13925_/Q vssd1 vssd1 vccd1 vccd1 hold2003/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09893_ _09995_/A _09892_/C _09892_/A vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2014 _07751_/X vssd1 vssd1 vccd1 vccd1 _14367_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _13934_/Q vssd1 vssd1 vccd1 vccd1 hold2025/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2036 _11955_/X vssd1 vssd1 vccd1 vccd1 _14775_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _07029_/X vssd1 vssd1 vccd1 vccd1 _13846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2047 _14735_/Q vssd1 vssd1 vccd1 vccd1 hold2047/X sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ _08526_/B _08842_/X _08843_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _08844_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1313 _15277_/Q vssd1 vssd1 vccd1 vccd1 hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _07088_/X vssd1 vssd1 vccd1 vccd1 _13901_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1324 _13692_/X vssd1 vssd1 vccd1 vccd1 _15398_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 _14216_/Q vssd1 vssd1 vccd1 vccd1 hold2069/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 _14671_/Q vssd1 vssd1 vccd1 vccd1 hold1335/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1346 _07775_/X vssd1 vssd1 vccd1 vccd1 _14391_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1357 _13804_/Q vssd1 vssd1 vccd1 vccd1 hold1357/X sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ _08776_/B _09858_/A _09858_/B _08776_/A vssd1 vssd1 vccd1 vccd1 _08775_/X
+ sky130_fd_sc_hd__a22o_1
Xhold1368 _07618_/X vssd1 vssd1 vccd1 vccd1 _14241_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout463_A _07045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1379 _14685_/Q vssd1 vssd1 vccd1 vccd1 hold1379/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ hold463/X _13732_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold464/A sky130_fd_sc_hd__mux2_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10655__A1 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10655__B2 _15207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_A _15202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ hold611/X _13729_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold612/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07520__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_A _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07588_ _13727_/A1 hold1049/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07588_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09327_ _09324_/X _09325_/Y _09186_/X _09190_/B vssd1 vssd1 vccd1 vccd1 _09328_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_193_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08076__A2 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _09255_/Y _09256_/X _09135_/X _09137_/X vssd1 vssd1 vccd1 vccd1 _09259_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08209_ _08209_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09025__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ _09186_/X _09187_/Y _09055_/B _09056_/Y vssd1 vssd1 vccd1 vccd1 _09190_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09025__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11220_ _11220_/A _11220_/B _11331_/B _11220_/D vssd1 vssd1 vccd1 vccd1 _11455_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_181_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07619__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _11577_/A _14967_/Q _10961_/X _10781_/B _14969_/Q vssd1 vssd1 vccd1 vccd1
+ _11156_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10102_ _11493_/A _10101_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _10102_/Y sky130_fd_sc_hd__o21ai_1
X_11082_ _11082_/A _11082_/B _11082_/C vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_41_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12332__A1 _13374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _10033_/A _10142_/A _11537_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _10141_/A
+ sky130_fd_sc_hd__nand4_1
X_14910_ _14971_/CLK _14910_/D vssd1 vssd1 vccd1 vccd1 _14910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2570 hold2858/X vssd1 vssd1 vccd1 vccd1 _07903_/C sky130_fd_sc_hd__clkbuf_2
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _14842_/CLK _14841_/D vssd1 vssd1 vccd1 vccd1 _14841_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2581 _07925_/X vssd1 vssd1 vccd1 vccd1 _07926_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2592 _12173_/X vssd1 vssd1 vccd1 vccd1 _14897_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1880 _07025_/X vssd1 vssd1 vccd1 vccd1 _13842_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _15450_/CLK _14772_/D vssd1 vssd1 vccd1 vccd1 _14772_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1891 _14589_/Q vssd1 vssd1 vccd1 vccd1 hold1891/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11984_ hold793/X _13673_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 hold794/A sky130_fd_sc_hd__mux2_1
XFILLER_0_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13723_ hold1047/X hold465/X _13732_/S vssd1 vssd1 vccd1 vccd1 _13723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _11493_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13091__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ hold1155/X _13654_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 _13654_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _10866_/A _10866_/B _10866_/C vssd1 vssd1 vccd1 vccd1 _10868_/A sky130_fd_sc_hd__and3_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _12327_/A _12604_/X _12602_/X vssd1 vssd1 vccd1 vccd1 _13151_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _10405_/B _13797_/A2 _13584_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15318_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ _11594_/A _11563_/A _11606_/B _11570_/B vssd1 vssd1 vccd1 vccd1 _10797_/X
+ sky130_fd_sc_hd__and4_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10447__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15324_/CLK _15324_/D vssd1 vssd1 vccd1 vccd1 _15324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ _12692_/A1 _12535_/X _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12536_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_164_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__D _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15255_ _15256_/CLK hold100/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12435__S _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ _12642_/A1 _12466_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12467_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10744__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12246__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12020__A0 hold2617/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07529__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14206_ _15434_/CLK _14206_/D vssd1 vssd1 vccd1 vccd1 _14206_/Q sky130_fd_sc_hd__dfxtp_1
X_11418_ _11418_/A _11551_/A _11418_/C vssd1 vssd1 vccd1 vccd1 _11551_/B sky130_fd_sc_hd__nand3_1
X_15186_ _15190_/CLK _15186_/D vssd1 vssd1 vccd1 vccd1 _15186_/Q sky130_fd_sc_hd__dfxtp_2
X_12398_ hold203/A hold403/A hold971/A _13961_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12398_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08775__B1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ _15456_/CLK _14137_/D vssd1 vssd1 vccd1 vccd1 _14137_/Q sky130_fd_sc_hd__dfxtp_1
X_11349_ _11620_/A _11614_/B _11188_/X _11189_/X _11564_/B vssd1 vssd1 vccd1 vccd1
+ _11354_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_120_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ _15225_/CLK _14068_/D vssd1 vssd1 vccd1 vccd1 _14068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ _13100_/S0 _13014_/X _13018_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _13020_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08560_ _14664_/Q _13937_/Q _15438_/Q _13905_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08561_/B sky130_fd_sc_hd__mux4_1
X_07511_ _07744_/A _14089_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__or3_2
X_08491_ _08491_/A _08491_/B _08491_/C vssd1 vssd1 vccd1 vccd1 _08492_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07442_ _08107_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14072_/D sky130_fd_sc_hd__and2_1
XFILLER_0_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ _15347_/Q _14060_/Q vssd1 vssd1 vccd1 vccd1 _07373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_175_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09112_ _10430_/B1 _09105_/Y _09107_/Y _09109_/Y _09111_/Y vssd1 vssd1 vccd1 vccd1
+ _09112_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_162_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09043_ _10185_/A _10022_/B _09043_/C _09167_/A vssd1 vssd1 vccd1 vccd1 _09167_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_161_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10654__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold410 hold410/A vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold432/A vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold443 hold443/A vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__buf_1
XANTENNA__12562__A1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10804__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold454 hold454/A vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold465 hold465/A vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold476 hold476/A vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 hold487/A vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 hold498/A vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ _11507_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09945_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout580_A _15219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11485__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _10115_/B _10033_/A _14956_/Q _14957_/Q vssd1 vssd1 vccd1 vccd1 _10030_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _07723_/X vssd1 vssd1 vccd1 vccd1 _14342_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07174__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1121 _14371_/Q vssd1 vssd1 vccd1 vccd1 hold1121/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 _07686_/X vssd1 vssd1 vccd1 vccd1 _14306_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _08717_/B _08717_/Y _08824_/X _08826_/Y vssd1 vssd1 vccd1 vccd1 _08829_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 _14215_/Q vssd1 vssd1 vccd1 vccd1 hold1143/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout845_A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 _07187_/X vssd1 vssd1 vccd1 vccd1 _13994_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 _15326_/Q vssd1 vssd1 vccd1 vccd1 _07422_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1176 _13653_/X vssd1 vssd1 vccd1 vccd1 _15360_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 _14485_/Q vssd1 vssd1 vccd1 vccd1 hold1187/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08981_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _08758_/X sky130_fd_sc_hd__or2_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _13475_/X vssd1 vssd1 vccd1 vccd1 _15234_/D sky130_fd_sc_hd__buf_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07709_ hold1219/X _13748_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 _07709_/X sky130_fd_sc_hd__mux2_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08689_/A _08689_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08691_/A sky130_fd_sc_hd__and3_1
XANTENNA__10829__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _10675_/Y _10676_/X _10719_/C _10719_/D vssd1 vssd1 vccd1 vccd1 _10720_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10666_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ _14807_/Q hold683/A _14647_/Q _14743_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _10583_/B sky130_fd_sc_hd__mux4_1
X_13370_ _13373_/A _13370_/B vssd1 vssd1 vccd1 vccd1 _15161_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _12317_/X _12318_/X _12320_/X _12319_/X _12669_/A1 _12700_/S1 vssd1 vssd1
+ vccd1 vccd1 _12321_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12228__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A0 _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ _15040_/CLK _15040_/D vssd1 vssd1 vccd1 vccd1 _15040_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_181_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12252_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12252_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08034__A _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10283__B _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11203_ _11588_/A _11537_/A _11623_/B _11409_/A vssd1 vssd1 vccd1 vccd1 _11206_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12553__B2 _13181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12183_ hold2555/X _12195_/A2 _12182_/X _13491_/A vssd1 vssd1 vccd1 vccd1 _12183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_61_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__A2 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13594__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _15419_/Q _14554_/Q hold513/A _14778_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11134_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07980__A1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ _11065_/A _11240_/A _11065_/C vssd1 vssd1 vccd1 vccd1 _11240_/B sky130_fd_sc_hd__nand3_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12856__A2 _13161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12400__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07084__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _10126_/B _11168_/A _11606_/A _10126_/A vssd1 vssd1 vccd1 vccd1 _10019_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_76_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output228_A _15459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _14840_/CLK _14824_/D vssd1 vssd1 vccd1 vccd1 _14824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _15394_/CLK _14755_/D vssd1 vssd1 vccd1 vccd1 _14755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08288__A2 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ hold1351/X _13656_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09485__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13706_ hold2157/X _13739_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__mux2_1
X_10918_ _10916_/Y _10917_/X _11640_/B1 _10915_/X vssd1 vssd1 vccd1 vccd1 _10918_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14686_ _14750_/CLK hold344/X vssd1 vssd1 vccd1 vccd1 hold343/A sky130_fd_sc_hd__dfxtp_1
X_11898_ _13653_/A1 hold2017/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_134_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ _08107_/A _13625_/C _13636_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15351_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _10848_/A _10848_/B _10848_/C vssd1 vssd1 vccd1 vccd1 _10850_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_14_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _14440_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13568_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08996__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12792__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ _15309_/CLK _15307_/D vssd1 vssd1 vccd1 vccd1 _15307_/Q sky130_fd_sc_hd__dfxtp_1
X_12519_ _12669_/A1 _12514_/X _12518_/X _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12520_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10474__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13499_ _13499_/A _13499_/B vssd1 vssd1 vccd1 vccd1 _13499_/X sky130_fd_sc_hd__and2_1
XFILLER_0_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_149_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ _15248_/CLK _15238_/D vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11289__B _13464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12544__A1 _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15169_ _15365_/CLK _15169_/D vssd1 vssd1 vccd1 vccd1 _15169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07991_ _08760_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _07991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09730_ _09731_/A _09731_/B vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__nand2b_1
X_06942_ _06942_/A vssd1 vssd1 vccd1 vccd1 _06942_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _09661_/A _11536_/B _09661_/C _09813_/A vssd1 vssd1 vccd1 vccd1 _09813_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13724__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08612_ _08612_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _08614_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09592_/X sky130_fd_sc_hd__or2_2
XFILLER_0_94_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07722__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08543_ _13570_/B _08541_/Y _08542_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _08543_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08474_ _08474_/A _08474_/B vssd1 vssd1 vccd1 vccd1 _08509_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_175_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _07425_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _07425_/X sky130_fd_sc_hd__and2_1
XFILLER_0_190_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12458__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _11894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07356_ _15340_/Q _15330_/Q _15339_/Q vssd1 vssd1 vccd1 vccd1 _07362_/D sky130_fd_sc_hd__or3b_1
XANTENNA__09876__C _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11130__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07287_ _07326_/A vssd1 vssd1 vccd1 vccd1 _07287_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07169__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _10166_/A _09026_/B _09858_/C _09709_/B vssd1 vssd1 vccd1 vccd1 _09027_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout795_A _14491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout720 _14965_/Q vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__buf_4
Xfanout731 _14958_/Q vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__buf_4
Xfanout742 _14954_/Q vssd1 vssd1 vccd1 vccd1 _10304_/D sky130_fd_sc_hd__clkbuf_4
X_09928_ _09919_/B _09773_/B _10744_/A vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12104__A _14992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout753 _14951_/Q vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__buf_4
Xfanout764 _14947_/Q vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__clkbuf_8
Xfanout775 _14945_/Q vssd1 vssd1 vccd1 vccd1 _11333_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout786 _14941_/Q vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09859_ _09709_/B _09858_/X _09857_/X vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__a21bo_1
Xfanout797 _14490_/Q vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__buf_8
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08062__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07714__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12870_/A _12870_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _12877_/B sky130_fd_sc_hd__or3b_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07632__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ hold919/X _13741_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold920/A sky130_fd_sc_hd__mux2_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _12284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_124 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12697__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ _15405_/CLK _14540_/D vssd1 vssd1 vccd1 vccd1 _14540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_168 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _13705_/A1 hold1411/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11752_/X sky130_fd_sc_hd__mux2_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10278__B _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10878_/B _10702_/C _10702_/A vssd1 vssd1 vccd1 vccd1 _10704_/C sky130_fd_sc_hd__a21o_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14471_ _15405_/CLK _14471_/D vssd1 vssd1 vccd1 vccd1 _14471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _13714_/A1 hold1393/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12449__S1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13422_ _13450_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13422_/Y sky130_fd_sc_hd__nand2_1
X_10634_ _10633_/B _10633_/C _10633_/A vssd1 vssd1 vccd1 vccd1 _10635_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13353_ _13360_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _15144_/D sky130_fd_sc_hd__nor2_1
X_10565_ _12256_/A _10563_/X _10564_/Y _12221_/B vssd1 vssd1 vccd1 vccd1 _10565_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _07439_/A hold277/A _06938_/Y _15350_/Q vssd1 vssd1 vccd1 vccd1 _12304_/X
+ sky130_fd_sc_hd__o22a_1
X_13284_ _13287_/A _13284_/B vssd1 vssd1 vccd1 vccd1 _15114_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10496_ _10496_/A _10496_/B _10482_/Y vssd1 vssd1 vccd1 vccd1 _10498_/B sky130_fd_sc_hd__nor3b_2
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output178_A _15189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15023_ _15188_/CLK _15023_/D vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
X_12235_ hold883/A _15262_/Q _15070_/Q _14363_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12235_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12621__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12166_ _14894_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__or2_1
X_11117_ _13750_/A _13370_/B _11116_/X vssd1 vssd1 vccd1 vccd1 _11117_/Y sky130_fd_sc_hd__o21ai_1
X_12097_ hold2398/X _12099_/A2 _12096_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12097_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12829__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ _11340_/A _15224_/Q vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__nand2_1
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09026__C _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 dmemresp_rdata[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07542__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ _15063_/CLK _14807_/D vssd1 vssd1 vccd1 vccd1 _14807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ hold1337/X hold775/X hold1687/X hold2235/X _12991_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12999_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_176_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09042__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _15378_/CLK hold866/X vssd1 vssd1 vccd1 vccd1 hold865/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08666__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14669_ _15445_/CLK _14669_/D vssd1 vssd1 vccd1 vccd1 _14669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07210_ hold775/X _13711_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold776/A sky130_fd_sc_hd__mux2_1
X_08190_ _08197_/A _08187_/X _08189_/X vssd1 vssd1 vccd1 vccd1 _08190_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07141_ _13742_/A1 hold1721/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07141_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09630__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15210__D _15210_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09630__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ hold2765/A hold2297/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput301 _14863_/Q vssd1 vssd1 vccd1 vccd1 out1[18] sky130_fd_sc_hd__buf_12
XANTENNA__12517__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput312 _14873_/Q vssd1 vssd1 vccd1 vccd1 out1[28] sky130_fd_sc_hd__buf_12
XFILLER_0_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13719__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput323 _14854_/Q vssd1 vssd1 vccd1 vccd1 out1[9] sky130_fd_sc_hd__buf_12
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput334 _14832_/Q vssd1 vssd1 vccd1 vccd1 out2[19] sky130_fd_sc_hd__buf_12
XFILLER_0_100_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput345 _14842_/Q vssd1 vssd1 vccd1 vccd1 out2[29] sky130_fd_sc_hd__buf_12
XFILLER_0_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07717__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08402__A _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07944__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07974_ _07974_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07975_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_199_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09713_ _09864_/A _09714_/C _09714_/D _09714_/A vssd1 vssd1 vccd1 vccd1 _09715_/B
+ sky130_fd_sc_hd__a22o_1
X_06925_ _09941_/A vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__inv_4
XFILLER_0_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13454__S _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_A _13502_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07960__B _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ hold805/A _14222_/Q hold515/A _14476_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09645_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09575_ _09434_/X _09436_/X _09573_/Y _09574_/X vssd1 vssd1 vccd1 vccd1 _09575_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout543_A _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08526_ _08526_/A _08526_/B vssd1 vssd1 vccd1 vccd1 _08526_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12453__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08457_ hold821/A _14212_/Q hold899/A _14466_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08458_/B sky130_fd_sc_hd__mux4_1
XANTENNA__08791__B _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout808_A _14489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07408_ _07408_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07408_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12205__B1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _09026_/B _09138_/A _08702_/B _08908_/A vssd1 vssd1 vccd1 vccd1 _08389_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10826__B _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11559__A2 _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07339_ hold573/A hold261/A _07855_/A vssd1 vssd1 vccd1 vccd1 _07849_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13202__B _13202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__A1 _11287_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11003__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10350_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ _09009_/A _09136_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _09011_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ _10282_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10463_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09385__B1 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ hold2617/X hold2682/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07627__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08312__A _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__A1 _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10090__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _10425_/S1 vssd1 vssd1 vccd1 vccd1 _10429_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout561 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _08763_/S0 sky130_fd_sc_hd__clkbuf_16
Xfanout572 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _11316_/S0 sky130_fd_sc_hd__clkbuf_8
Xfanout583 _10338_/C vssd1 vssd1 vccd1 vccd1 _11564_/B sky130_fd_sc_hd__clkbuf_8
X_13971_ _14602_/CLK _13971_/D vssd1 vssd1 vccd1 vccd1 _13971_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout594 _15213_/Q vssd1 vssd1 vccd1 vccd1 _09979_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__12141__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A2 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _14805_/Q _14517_/Q hold919/A _14741_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12922_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12692__B1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08685__C _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12853_ _13705_/A1 _13103_/A2 _13078_/B1 _13193_/B vssd1 vssd1 vccd1 vccd1 _12853_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ hold1515/X _13691_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11804_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13641__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12784_ hold511/X _13913_/Q _12791_/S vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__mux2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _15196_/CLK hold876/X vssd1 vssd1 vccd1 vccd1 hold875/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _13721_/A1 hold2195/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11735_/X sky130_fd_sc_hd__mux2_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ _15324_/CLK _14454_/D vssd1 vssd1 vccd1 vccd1 _14454_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _13730_/A1 hold1069/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11666_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _13479_/A _13405_/B vssd1 vssd1 vccd1 vccd1 _15196_/D sky130_fd_sc_hd__and2_1
X_10617_ _11573_/A _11594_/A _11606_/B _11570_/B vssd1 vssd1 vccd1 vccd1 _10619_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_25_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14385_ _15408_/CLK _14385_/D vssd1 vssd1 vccd1 vccd1 _14385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12009__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11597_ _11597_/A _14968_/Q vssd1 vssd1 vccd1 vccd1 _11599_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15030__D _15030_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ input153/X fanout5/X fanout3/X input121/X vssd1 vssd1 vccd1 vccd1 _13336_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10222__A2 _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ _10548_/A _10548_/B _10548_/C _10548_/D vssd1 vssd1 vccd1 vccd1 _10548_/X
+ sky130_fd_sc_hd__or4_2
Xclkbuf_4_5__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13267_ input159/X fanout6/X fanout4/X input127/X vssd1 vssd1 vccd1 vccd1 _13267_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10479_ _10303_/X _10305_/X _10477_/Y _10478_/X vssd1 vssd1 vccd1 vccd1 _10479_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15006_ _15268_/CLK _15006_/D vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07537__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _12241_/A _12218_/B vssd1 vssd1 vccd1 vccd1 _12219_/D sky130_fd_sc_hd__nand2_1
XANTENNA__11567__B _15228_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__B _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _13404_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _15063_/D sky130_fd_sc_hd__and2_1
XFILLER_0_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ hold2602/X _12173_/A2 _12148_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12149_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1709 _14373_/Q vssd1 vssd1 vccd1 vccd1 hold1709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07690_ hold365/X _13663_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold366/A sky130_fd_sc_hd__mux2_1
XFILLER_0_189_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09360_ _10426_/A _09359_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08892__A _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _08310_/A _08310_/B _08310_/C vssd1 vssd1 vccd1 vccd1 _08312_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12986__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09291_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08242_ _08243_/B _08242_/B vssd1 vssd1 vccd1 vccd1 _08242_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_129_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_24 _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_35 _14928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__B _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_46 _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07301__A _15219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 _07326_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _12221_/B _08244_/C _08172_/X _08526_/B hold2761/X vssd1 vssd1 vccd1 vccd1
+ _08173_/X sky130_fd_sc_hd__a32o_1
XANTENNA_68 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_79 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12833__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1_N _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _13725_/A1 hold2025/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07124_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07055_ _13512_/A0 hold1839/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07055_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12353__S _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12597__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput164 _15176_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[11] sky130_fd_sc_hd__buf_12
XANTENNA__07917__A1 _07431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput175 _15186_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[21] sky130_fd_sc_hd__buf_12
XANTENNA_fanout493_A _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 _15196_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[31] sky130_fd_sc_hd__buf_12
XFILLER_0_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput197 _14180_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[10] sky130_fd_sc_hd__buf_12
X_07957_ _07958_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__or2_1
XFILLER_0_199_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout758_A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__C1 _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _15345_/Q vssd1 vssd1 vccd1 vccd1 _06908_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_97_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07888_ _08677_/A _11566_/A _07889_/C vssd1 vssd1 vccd1 vccd1 _07890_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08342__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09627_ _09775_/A _09775_/B _09490_/Y vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_210_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09558_ _09557_/B _09557_/C _09557_/A vssd1 vssd1 vccd1 vccd1 _09558_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08509_ _08509_/A _08509_/B vssd1 vssd1 vccd1 vccd1 _08511_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12431__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12521__S0 _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ _09218_/A _09349_/A _09488_/Y vssd1 vssd1 vccd1 vccd1 _09491_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11520_ _11467_/A _11466_/B _11466_/A vssd1 vssd1 vccd1 vccd1 _11521_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout3_A fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _11183_/A _11183_/Y _11607_/B _11450_/X vssd1 vssd1 vccd1 vccd1 _11453_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_0_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08026__B _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10275__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__S1 _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07605__A0 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _10228_/B _09927_/B _09919_/B _09773_/B _10744_/A vssd1 vssd1 vccd1 vccd1
+ _10402_/X sky130_fd_sc_hd__o41a_1
X_14170_ _15268_/CLK hold174/X vssd1 vssd1 vccd1 vccd1 _14170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ _11382_/A _11382_/B vssd1 vssd1 vccd1 vccd1 _11383_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13121_ _13490_/A hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__and2_1
X_10333_ _10333_/A _10333_/B _10333_/C vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_103_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09138__A _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _13102_/A _13052_/B _13052_/C vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__and3_1
X_10264_ _09763_/A _09763_/B _10071_/X _10265_/B vssd1 vssd1 vccd1 vccd1 _10268_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11165__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A _14428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12003_ _12063_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _14814_/D sky130_fd_sc_hd__and2_1
XANTENNA__08030__B1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10195_ _09987_/Y _09989_/X _10193_/Y _10194_/X vssd1 vssd1 vccd1 vccd1 _10198_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_108_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08696__B _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13457__A2 _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout380 _12309_/Y vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_13__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_76_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout391 _07900_/B vssd1 vssd1 vccd1 vccd1 _11288_/A1 sky130_fd_sc_hd__buf_12
XFILLER_0_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13954_ _15455_/CLK _13954_/D vssd1 vssd1 vccd1 vccd1 _13954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07092__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ _13080_/A1 _12904_/X _12902_/X vssd1 vssd1 vccd1 vccd1 _13163_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13885_ _15408_/CLK _13885_/D vssd1 vssd1 vccd1 vccd1 _13885_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08884__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12445__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ _12917_/A1 _12835_/X _12844_/A1 vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12417__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13614__C1 _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12767_ _12917_/A1 _12766_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12767_/X sky130_fd_sc_hd__a21o_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10979__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08192__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ _15369_/CLK hold726/X vssd1 vssd1 vccd1 vccd1 hold725/A sky130_fd_sc_hd__dfxtp_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11718_ hold1483/X _13738_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 _11718_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12698_ hold249/A _14313_/Q _14604_/Q _13973_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12698_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12595__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14437_ _15309_/CLK _14437_/D vssd1 vssd1 vccd1 vccd1 _14437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ _10233_/A _11643_/Y _11648_/X _11491_/X vssd1 vssd1 vccd1 vccd1 _11649_/X
+ sky130_fd_sc_hd__a31o_1
Xinput11 dmemresp_rdata[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput22 dmemresp_rdata[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 imemresp_data[0] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 imemresp_data[1] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput55 imemresp_data[2] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
X_14368_ _15364_/CLK _14368_/D vssd1 vssd1 vccd1 vccd1 _14368_/Q sky130_fd_sc_hd__dfxtp_1
Xinput66 in0[10] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_1
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput77 in0[20] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold806 hold806/A vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold817 hold817/A vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 in0[30] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_1
X_13319_ input82/X fanout2/X _13318_/X vssd1 vssd1 vccd1 vccd1 _13320_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11578__A _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold828 hold828/A vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 in1[11] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
Xhold839 hold839/A vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _15364_/CLK hold744/X vssd1 vssd1 vccd1 vccd1 hold743/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11297__B _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2207 _13938_/Q vssd1 vssd1 vccd1 vccd1 hold2207/X sky130_fd_sc_hd__dlygate4sd3_1
X_08860_ _11104_/A _12273_/B _08859_/X vssd1 vssd1 vccd1 vccd1 _08860_/X sky130_fd_sc_hd__a21bo_1
Xhold2218 _06980_/X vssd1 vssd1 vccd1 vccd1 _13799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2229 _13944_/Q vssd1 vssd1 vccd1 vccd1 hold2229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07811_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__nor2_4
Xhold1506 _11785_/X vssd1 vssd1 vccd1 vccd1 _14610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 _14238_/Q vssd1 vssd1 vccd1 vccd1 hold1517/X sky130_fd_sc_hd__dlygate4sd3_1
X_08791_ _09661_/A _09858_/C vssd1 vssd1 vccd1 vccd1 _08794_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1528 _07490_/X vssd1 vssd1 vccd1 vccd1 _14118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _14702_/Q vssd1 vssd1 vccd1 vccd1 hold1539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07742_ hold1463/X _13748_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07742_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12656__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07673_ hold599/X _13745_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 hold600/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_185_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15365_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09412_ _09411_/B _09411_/C _09411_/A vssd1 vssd1 vccd1 vccd1 _09412_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13732__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07730__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _11288_/A1 _09342_/X _09245_/X vssd1 vssd1 vccd1 vccd1 _12277_/B sky130_fd_sc_hd__a21o_4
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13081__B1 _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12348__S _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09274_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__and2_1
XFILLER_0_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08127__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08225_ _08226_/A _08226_/B _08226_/C vssd1 vssd1 vccd1 vccd1 _08225_/X sky130_fd_sc_hd__and3_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout506_A _06926_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08156_ _08156_/A _08156_/B _08209_/B vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__and3_1
XFILLER_0_209_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07107_ _13743_/A1 hold2211/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07107_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08260__B1 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08087_ _10873_/A _09138_/A _08161_/A _08088_/D vssd1 vssd1 vccd1 vccd1 _08089_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07177__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ hold739/X _11921_/A0 _07044_/S vssd1 vssd1 vccd1 vccd1 hold740/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout875_A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11698__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2730 _12454_/X vssd1 vssd1 vccd1 vccd1 hold2730/X sky130_fd_sc_hd__buf_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2741 _15188_/Q vssd1 vssd1 vccd1 vccd1 hold2741/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2752 _10918_/X vssd1 vssd1 vccd1 vccd1 _13401_/B sky130_fd_sc_hd__buf_1
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08989_/Y sky130_fd_sc_hd__nor2_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2763 _15186_/Q vssd1 vssd1 vccd1 vccd1 hold2763/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2774 _14491_/Q vssd1 vssd1 vccd1 vccd1 hold2774/X sky130_fd_sc_hd__clkbuf_2
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2785 _11641_/X vssd1 vssd1 vccd1 vccd1 _13405_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2796 _15126_/Q vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12112__A _12112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _10951_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10952_/B sky130_fd_sc_hd__or2_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11373__D _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_176_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_211_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11870__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ hold695/X _13736_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold696/A sky130_fd_sc_hd__mux2_1
XFILLER_0_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10882_ _11517_/A _11586_/B _10881_/C _10881_/D vssd1 vssd1 vccd1 vccd1 _10882_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_74_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07640__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _15370_/Q _15273_/Q _15081_/Q _14374_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12621_/X sky130_fd_sc_hd__mux4_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12258__S _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15340_ _15340_/CLK _15340_/D vssd1 vssd1 vccd1 vccd1 _15340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__A1 _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ _13027_/A _12552_/B _12552_/C vssd1 vssd1 vccd1 vccd1 _12552_/X sky130_fd_sc_hd__and3_1
XANTENNA__10286__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11503_ _13893_/Q _14021_/Q hold871/A _13829_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11504_/B sky130_fd_sc_hd__mux4_1
X_15271_ _15416_/CLK _15271_/D vssd1 vssd1 vccd1 vccd1 _15271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12483_ hold519/A hold901/A hold543/A _14756_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12483_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14222_ _15410_/CLK _14222_/D vssd1 vssd1 vccd1 vccd1 _14222_/Q sky130_fd_sc_hd__dfxtp_1
X_11434_ _11434_/A _11575_/A _11434_/C vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__and3_1
XFILLER_0_110_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14153_ _15405_/CLK hold606/X vssd1 vssd1 vccd1 vccd1 hold605/A sky130_fd_sc_hd__dfxtp_1
X_11365_ _11365_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_100_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15243_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07087__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13104_ _11641_/X _13104_/A2 _13103_/X vssd1 vssd1 vccd1 vccd1 _13104_/X sky130_fd_sc_hd__a21o_1
X_10316_ _11569_/A _10316_/B _10483_/A _10316_/D vssd1 vssd1 vccd1 vccd1 _10483_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_131_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14084_ _14105_/CLK _14084_/D vssd1 vssd1 vccd1 vccd1 _14084_/Q sky130_fd_sc_hd__dfxtp_1
X_11296_ _13594_/A _11295_/B _07390_/A vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_output258_A _14432_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ hold877/A _13955_/Q _13041_/S vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__mux2_1
X_10247_ _14354_/Q _14258_/Q hold897/A _14130_/Q _10425_/S0 _10425_/S1 vssd1 vssd1
+ vccd1 vccd1 _10248_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12886__B1 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10178_ _10351_/A _15220_/Q vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_206_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14986_ _15243_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _14986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12733__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_167_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15276_/CLK sky130_fd_sc_hd__clkbuf_16
X_13937_ _15438_/CLK _13937_/D vssd1 vssd1 vccd1 vccd1 _13937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13868_ _15394_/CLK _13868_/D vssd1 vssd1 vccd1 vccd1 _13868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11580__B _14972_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _12844_/A1 _12814_/X _12818_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12820_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10477__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09806__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ _15261_/CLK _13799_/D vssd1 vssd1 vccd1 vccd1 _13799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ _08010_/A _08010_/B _08010_/C vssd1 vssd1 vccd1 vccd1 _08012_/C sky130_fd_sc_hd__nand3_1
XANTENNA__11800__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__B1 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2540_A _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 hold603/A vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold614 hold614/A vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold625 hold625/A vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 hold636/A vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10643__C _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 hold647/A vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold658 hold658/A vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _11335_/A _10338_/C _09959_/Y _10170_/A vssd1 vssd1 vccd1 vccd1 _09963_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_111_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold669 hold669/A vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08912_ _08912_/A _08912_/B _08912_/C vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__and3_1
XANTENNA__13727__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _09892_/A _09995_/A _09892_/C vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__and3_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2004 _07112_/X vssd1 vssd1 vccd1 vccd1 _13925_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 _15381_/Q vssd1 vssd1 vccd1 vccd1 hold2015/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07725__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2026 _07124_/X vssd1 vssd1 vccd1 vccd1 _13934_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08843_ _08843_/A _12256_/A vssd1 vssd1 vccd1 vccd1 _08843_/X sky130_fd_sc_hd__or2_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12972__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2037 _13990_/Q vssd1 vssd1 vccd1 vccd1 hold2037/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2048 _11914_/X vssd1 vssd1 vccd1 vccd1 _14735_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1303 _14662_/Q vssd1 vssd1 vccd1 vccd1 hold1303/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _13519_/X vssd1 vssd1 vccd1 vccd1 _15277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2059 _13907_/Q vssd1 vssd1 vccd1 vccd1 hold2059/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 _14396_/Q vssd1 vssd1 vccd1 vccd1 hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1336 _11848_/X vssd1 vssd1 vccd1 vccd1 _14671_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _09435_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _08778_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1347 _14344_/Q vssd1 vssd1 vccd1 vccd1 hold1347/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1358 _06985_/X vssd1 vssd1 vccd1 vccd1 _13804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1369 _14353_/Q vssd1 vssd1 vccd1 vccd1 hold1369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12724__S0 _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07725_ hold1347/X _13698_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 _07725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_158_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15432_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10104__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A2 _13387_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout456_A _07012_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13462__S _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10655__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ hold993/X _13728_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold994/A sky130_fd_sc_hd__mux2_1
XFILLER_0_192_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout623_A _15204_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07587_ _13693_/A1 hold577/X _07593_/S vssd1 vssd1 vccd1 vccd1 hold578/A sky130_fd_sc_hd__mux2_1
X_09326_ _09186_/X _09190_/B _09324_/X _09325_/Y vssd1 vssd1 vccd1 vccd1 _09328_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09257_ _09135_/X _09137_/X _09255_/Y _09256_/X vssd1 vssd1 vccd1 vccd1 _09257_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11710__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08208_ _13724_/A1 _12260_/A2 _12259_/A1 _13179_/B _08206_/Y vssd1 vssd1 vccd1 vccd1
+ _08208_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09025__A2 _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09188_ _09055_/B _09056_/Y _09186_/X _09187_/Y vssd1 vssd1 vccd1 vccd1 _09190_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_161_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08459__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08139_ _08139_/A _08214_/A vssd1 vssd1 vccd1 vccd1 _08156_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _11150_/A _11150_/B vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ hold679/A _14548_/Q hold325/A _14772_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10101_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ _11081_/A _11081_/B vssd1 vssd1 vccd1 vccd1 _11082_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__10850__A _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12541__S _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _11573_/A _14956_/Q _14957_/Q _10033_/A vssd1 vssd1 vccd1 vccd1 _10035_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2560 hold2856/X vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _14840_/CLK _14840_/D vssd1 vssd1 vccd1 vccd1 _14840_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2571 _15316_/Q vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2582 _07927_/Y vssd1 vssd1 vccd1 vccd1 _14426_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2593 _14992_/Q vssd1 vssd1 vccd1 vccd1 hold2593/X sky130_fd_sc_hd__buf_2
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1870 _07076_/X vssd1 vssd1 vccd1 vccd1 _13892_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1881 _14753_/Q vssd1 vssd1 vccd1 vccd1 hold1881/X sky130_fd_sc_hd__dlygate4sd3_1
X_14771_ _15449_/CLK _14771_/D vssd1 vssd1 vccd1 vccd1 _14771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11983_ hold1577/X _13705_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11983_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_149_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15079_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12777__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1892 _11764_/X vssd1 vssd1 vccd1 vccd1 _14589_/D sky130_fd_sc_hd__dlygate4sd3_1
X_13722_ hold661/X hold2783/X _13732_/S vssd1 vssd1 vccd1 vccd1 hold662/A sky130_fd_sc_hd__mux2_1
XFILLER_0_168_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10934_ hold371/A hold349/A hold363/A _14745_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _10935_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_169_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08466__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09151__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13653_ hold1175/X _13653_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 _13653_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_195_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10297__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10865_ _10681_/B _10681_/C _10681_/A vssd1 vssd1 vccd1 vccd1 _10866_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _13385_/B _12325_/B _12603_/X vssd1 vssd1 vccd1 vccd1 _12604_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13584_ _13584_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__or2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _11563_/A _11606_/B _11570_/B _11594_/A vssd1 vssd1 vccd1 vccd1 _10801_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15324_/CLK _15323_/D vssd1 vssd1 vccd1 vccd1 _15323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10447__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12535_ _14662_/Q _13935_/Q _12560_/S vssd1 vssd1 vccd1 vccd1 _12535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12716__S _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13401__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ _15254_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12466_ hold337/A hold913/A _12466_/S vssd1 vssd1 vccd1 vccd1 _12466_/X sky130_fd_sc_hd__mux2_1
X_14205_ _14397_/CLK _14205_/D vssd1 vssd1 vccd1 vccd1 _14205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11417_ _11416_/A _11608_/B _11416_/C vssd1 vssd1 vccd1 vccd1 _11418_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15185_ _15190_/CLK _15185_/D vssd1 vssd1 vccd1 vccd1 _15185_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12397_ _14784_/Q hold939/A hold923/A _14720_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12397_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08775__A1 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B2 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14136_ _14972_/CLK _14136_/D vssd1 vssd1 vccd1 vccd1 _14136_/Q sky130_fd_sc_hd__dfxtp_1
X_11348_ _11348_/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11356_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14067_ _15222_/CLK _14067_/D vssd1 vssd1 vccd1 vccd1 _14067_/Q sky130_fd_sc_hd__dfxtp_1
X_11279_ _11280_/B vssd1 vssd1 vccd1 vccd1 _11279_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13018_ _13099_/S1 _13015_/X _13017_/X vssd1 vssd1 vccd1 vccd1 _13018_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14969_ _14972_/CLK _14969_/D vssd1 vssd1 vccd1 vccd1 _14969_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_18_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07510_ _14088_/Q _11729_/B _14090_/Q vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__and3_2
XFILLER_0_57_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08490_ _08491_/A _08491_/B _08491_/C vssd1 vssd1 vccd1 vccd1 _08492_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ _12294_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14071_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13036__B1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10000__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07372_ _15347_/Q _14060_/Q vssd1 vssd1 vccd1 vccd1 _07372_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09111_ _09941_/A _09110_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09111_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10935__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13311__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ _10183_/A _09979_/B _09864_/A _10022_/A vssd1 vssd1 vccd1 vccd1 _09167_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__10270__B1 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10654__B _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold400 hold400/A vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold411 hold411/A vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold422/A vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold433 hold433/A vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold444 hold444/A vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold455 hold455/A vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/A vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold477 hold477/A vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ hold931/A hold699/A hold501/A _14128_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _09945_/B sky130_fd_sc_hd__mux4_1
Xhold488 hold488/A vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09236__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _10033_/A _09724_/C _09724_/D _10115_/B vssd1 vssd1 vccd1 vccd1 _09878_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08140__A _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 _11837_/X vssd1 vssd1 vccd1 vccd1 _14660_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout573_A _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _14799_/Q vssd1 vssd1 vccd1 vccd1 hold1111/X sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ _08825_/B _08825_/C _08825_/A vssd1 vssd1 vccd1 vccd1 _08826_/Y sky130_fd_sc_hd__a21oi_2
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _07755_/X vssd1 vssd1 vccd1 vccd1 _14371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _15440_/Q vssd1 vssd1 vccd1 vccd1 hold1133/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 _07591_/X vssd1 vssd1 vccd1 vccd1 _14215_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 _15361_/Q vssd1 vssd1 vccd1 vccd1 hold1155/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1166 _07422_/X vssd1 vssd1 vccd1 vccd1 _14052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ hold785/A hold725/A _14634_/Q _14730_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08758_/B sky130_fd_sc_hd__mux4_1
Xhold1177 _13985_/Q vssd1 vssd1 vccd1 vccd1 hold1177/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1188 _11682_/X vssd1 vssd1 vccd1 vccd1 _14485_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1199 _13875_/Q vssd1 vssd1 vccd1 vccd1 hold1199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11705__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07708_ hold1229/X _13681_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 _07708_/X sky130_fd_sc_hd__mux2_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08586_/A _08586_/B _08586_/C vssd1 vssd1 vccd1 vccd1 _08689_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__08286__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10829__B _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07639_ hold667/X _13745_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold668/A sky130_fd_sc_hd__mux2_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ _10648_/X _10650_/B vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_193_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09309_ _09175_/B _09178_/B _09307_/X _09308_/Y vssd1 vssd1 vccd1 vccd1 _09309_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12250__A1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ hold315/A hold449/A hold523/A _14388_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _10581_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09651__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _13862_/Q _13990_/Q _13830_/Q _13798_/Q _12365_/S0 _12365_/S1 vssd1 vssd1
+ vccd1 vccd1 _12320_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_180_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10564__B _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ _12234_/X _12241_/Y _12250_/X _12241_/A vssd1 vssd1 vccd1 vccd1 _12252_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10239__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10283__C _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ _11407_/A _11588_/B _10979_/X _10980_/X _11606_/B vssd1 vssd1 vccd1 vccd1
+ _11207_/A sky130_fd_sc_hd__a32o_1
XANTENNA__12553__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ _14902_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _11504_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11133_/Y sky130_fd_sc_hd__nor2_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ _11063_/B _11242_/B _11063_/A vssd1 vssd1 vccd1 vccd1 _11065_/C sky130_fd_sc_hd__a21o_1
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09801__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__xnor2_2
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08985__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2390 hold2845/X vssd1 vssd1 vccd1 vccd1 _06904_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_203_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _14840_/CLK _14823_/D vssd1 vssd1 vccd1 vccd1 _14823_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08368__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11966_ hold1575/X _13655_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11966_/X sky130_fd_sc_hd__mux2_1
X_14754_ _14754_/CLK _14754_/D vssd1 vssd1 vccd1 vccd1 _14754_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09485__A2 _13392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ _10951_/A _07296_/B _10602_/X _11640_/B1 vssd1 vssd1 vccd1 vccd1 _10917_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07496__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13705_ hold1813/X _13705_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13705_/X sky130_fd_sc_hd__mux2_1
X_14685_ _15426_/CLK _14685_/D vssd1 vssd1 vccd1 vccd1 _14685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11897_ _13652_/A1 hold2197/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13636_ input50/X _13636_/B vssd1 vssd1 vccd1 vccd1 _13636_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10848_ _10848_/A _10848_/B _10848_/C vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08445__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ _09083_/A _09222_/B _13566_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10779_ _11578_/A _14967_/Q _14968_/Q _11580_/A vssd1 vssd1 vccd1 vccd1 _10782_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08996__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ _12368_/A _12515_/X _12517_/X vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__a21o_1
X_15306_ _15309_/CLK _15306_/D vssd1 vssd1 vccd1 vccd1 _15306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13498_ _13499_/A hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__and2_1
XANTENNA__10474__B _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ _13867_/Q hold387/A _13835_/Q _13803_/Q _12460_/S _12689_/S1 vssd1 vssd1
+ vccd1 vccd1 _12449_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_48_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15237_ _15246_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15168_ _15365_/CLK _15168_/D vssd1 vssd1 vccd1 vccd1 _15168_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11752__A0 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ _14602_/CLK _14119_/D vssd1 vssd1 vccd1 vccd1 _14119_/Q sky130_fd_sc_hd__dfxtp_1
X_07990_ _08201_/A _07987_/X _07989_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _07991_/B
+ sky130_fd_sc_hd__o211a_1
X_15099_ _15457_/CLK hold452/X vssd1 vssd1 vccd1 vccd1 hold451/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06941_ _06941_/A vssd1 vssd1 vccd1 vccd1 _06941_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _09661_/A _11536_/B _09661_/C _09813_/A vssd1 vssd1 vccd1 vccd1 _09663_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08611_ _08612_/A _08612_/B vssd1 vssd1 vccd1 vccd1 _08611_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09591_ _09591_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09593_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _08542_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _08542_/X sky130_fd_sc_hd__or2_1
XANTENNA__12210__A _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08133__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07304__A _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _08473_/A _08473_/B _08503_/B vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__or3b_1
XANTENNA__12480__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__B1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13740__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _07424_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _14054_/D sky130_fd_sc_hd__and2_1
XFILLER_0_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07355_ _08635_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07355_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09876__D _14957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A _13650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07286_ _15228_/Q _14972_/Q vssd1 vssd1 vccd1 vccd1 _07326_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09025_ _09026_/B _09858_/C _09709_/B _08908_/A vssd1 vssd1 vccd1 vccd1 _09027_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08739__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13732__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__buf_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout710 _13721_/A1 vssd1 vssd1 vccd1 vccd1 _13655_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout721 _14964_/Q vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__07185__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 _11623_/B vssd1 vssd1 vccd1 vccd1 _09724_/D sky130_fd_sc_hd__buf_4
X_09927_ _10744_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _10401_/A sky130_fd_sc_hd__xnor2_1
Xfanout743 _14953_/Q vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__buf_4
Xfanout754 _14950_/Q vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__buf_4
XANTENNA__12104__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 _09542_/A vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__clkbuf_8
Xfanout776 _14944_/Q vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__clkbuf_8
X_09858_ _09858_/A _09858_/B _09858_/C vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__and3_1
Xfanout787 _14941_/Q vssd1 vssd1 vccd1 vccd1 _11567_/A sky130_fd_sc_hd__clkbuf_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 _06943_/A vssd1 vssd1 vccd1 vccd1 _12917_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_198_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _09571_/A _08809_/B _09714_/A _08809_/D vssd1 vssd1 vccd1 vccd1 _08922_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _10244_/A _09786_/X _09788_/X vssd1 vssd1 vccd1 vccd1 _09789_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_103 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ hold847/X _13674_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold848/A sky130_fd_sc_hd__mux2_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _12284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__A _12120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_125 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_136 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ _13704_/A1 hold1461/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__mux2_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _14776_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10702_ _10702_/A _10878_/B _10702_/C vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__nand3_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _15436_/CLK _14470_/D vssd1 vssd1 vccd1 vccd1 _14470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11682_ _13746_/A1 hold1187/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09219__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _08253_/B _13440_/S _13420_/Y _13178_/A vssd1 vssd1 vccd1 vccd1 _15204_/D
+ sky130_fd_sc_hd__o211a_1
X_10633_ _10633_/A _10633_/B _10633_/C vssd1 vssd1 vccd1 vccd1 _10819_/A sky130_fd_sc_hd__and3_1
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10234__B1 _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08978__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13352_ _13360_/A _13352_/B vssd1 vssd1 vccd1 vccd1 _15143_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ _10564_/A _11283_/S vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10785__A1 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12303_ _07438_/A _14032_/Q hold278/A _15348_/Q _12302_/X vssd1 vssd1 vccd1 vccd1
+ _12303_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_180_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13283_ input69/X fanout1/X _13282_/X vssd1 vssd1 vccd1 vccd1 _13284_/B sky130_fd_sc_hd__a21oi_1
X_10495_ _10494_/A _10494_/B _10494_/C vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__a21oi_1
X_15022_ _15278_/CLK _15022_/D vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__dfxtp_1
X_12234_ _12243_/A _12231_/Y _12233_/Y _06926_/A _12229_/Y vssd1 vssd1 vccd1 vccd1
+ _12234_/X sky130_fd_sc_hd__a311o_1
XANTENNA__11734__A0 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ hold2471/X _12173_/A2 _12164_/X _13129_/A vssd1 vssd1 vccd1 vccd1 _12165_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07095__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11116_ _10233_/A _11295_/B _11114_/Y _11115_/Y vssd1 vssd1 vccd1 vccd1 _11116_/X
+ sky130_fd_sc_hd__o31a_1
X_12096_ _14988_/Q _12096_/B _12096_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12096_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _11047_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__or2_1
XFILLER_0_127_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09026__D _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__A1 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 dmemresp_rdata[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _15242_/CLK hold300/X vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ hold157/X hold1883/X hold623/X hold1177/X _12991_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12998_/X sky130_fd_sc_hd__mux4_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09042__C _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14737_ _15378_/CLK _14737_/D vssd1 vssd1 vccd1 vccd1 _14737_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12462__A1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _13704_/A1 hold1173/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_71_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _14972_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08761__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14668_ _15439_/CLK _14668_/D vssd1 vssd1 vccd1 vccd1 _14668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13619_ input35/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13619_/X sky130_fd_sc_hd__or2_1
XANTENNA__10485__A _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ _15400_/CLK _14599_/D vssd1 vssd1 vccd1 vccd1 _14599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07140_ _13741_/A1 hold1677/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07140_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09630__A2 _13444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ _11921_/A0 hold2255/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07071_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput302 _14864_/Q vssd1 vssd1 vccd1 vccd1 out1[19] sky130_fd_sc_hd__buf_12
Xoutput313 _14874_/Q vssd1 vssd1 vccd1 vccd1 out1[29] sky130_fd_sc_hd__buf_12
Xoutput324 _14813_/Q vssd1 vssd1 vccd1 vccd1 out2[0] sky130_fd_sc_hd__buf_12
XFILLER_0_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput335 _14814_/Q vssd1 vssd1 vccd1 vccd1 out2[1] sky130_fd_sc_hd__buf_12
XFILLER_0_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput346 _14815_/Q vssd1 vssd1 vccd1 vccd1 out2[2] sky130_fd_sc_hd__buf_12
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08402__B _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07973_ _07974_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__or2_1
X_09712_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09715_/A sky130_fd_sc_hd__and2_1
XANTENNA__13735__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11489__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06924_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__inv_2
XANTENNA__07157__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07733__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09643_ _10244_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09643_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09514__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout369_A _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09574_ _09864_/A _09712_/B _09573_/C _09573_/D vssd1 vssd1 vccd1 vccd1 _09574_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_180_clk_A clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08525_ _08521_/X _08523_/Y _08571_/B _10397_/A vssd1 vssd1 vccd1 vccd1 _08525_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout536_A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__B2 _13177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_A clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14844_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08752__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08456_ _12243_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08456_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_175_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07407_ _07407_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07407_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11008__A2 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12205__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _08908_/A _09026_/B _09138_/A _08702_/B vssd1 vssd1 vccd1 vccd1 _08389_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__10826__C _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07338_ _07903_/C _09344_/B _07336_/Y vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__A2 _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11003__B _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ _11537_/B _09724_/D vssd1 vssd1 vccd1 vccd1 _07271_/A sky130_fd_sc_hd__or2_1
XFILLER_0_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09008_ _09008_/A _09136_/A _09714_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09008_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13705__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10282_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09385__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12913__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08312__B _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_133_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _08763_/S1 vssd1 vssd1 vccd1 vccd1 _08990_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout551 _15423_/Q vssd1 vssd1 vccd1 vccd1 _10425_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout562 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _12237_/S sky130_fd_sc_hd__buf_8
X_13970_ _15432_/CLK _13970_/D vssd1 vssd1 vccd1 vccd1 _13970_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout573 _11501_/S0 vssd1 vssd1 vccd1 vccd1 _10930_/S0 sky130_fd_sc_hd__buf_8
Xfanout584 _15217_/Q vssd1 vssd1 vccd1 vccd1 _10338_/C sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_13_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 _09979_/C vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__clkbuf_8
X_12921_ hold843/A hold625/A hold741/A _14386_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12921_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12692__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08685__D _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_148_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12852_ _13102_/A _12852_/B _12852_/C vssd1 vssd1 vccd1 vccd1 _12852_/X sky130_fd_sc_hd__and3_1
XFILLER_0_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11803_ hold995/X _13657_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold996/A sky130_fd_sc_hd__mux2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ hold879/A _14544_/Q _14704_/Q _14768_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12783_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12444__A1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_28_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15351_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _13687_/A1 hold2163/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11734_/X sky130_fd_sc_hd__mux2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _15387_/CLK hold414/X vssd1 vssd1 vccd1 vccd1 hold413/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _13729_/A1 hold1803/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11665_/X sky130_fd_sc_hd__mux2_1
X_14453_ _15296_/CLK _14453_/D vssd1 vssd1 vccd1 vccd1 _14453_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_154_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ _11594_/A _11606_/B _11570_/B _11573_/A vssd1 vssd1 vccd1 vccd1 _10619_/C
+ sky130_fd_sc_hd__a22o_1
X_13404_ _13404_/A _13404_/B vssd1 vssd1 vccd1 vccd1 _15195_/D sky130_fd_sc_hd__and2_1
XFILLER_0_25_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14384_ _15441_/CLK _14384_/D vssd1 vssd1 vccd1 vccd1 _14384_/Q sky130_fd_sc_hd__dfxtp_1
X_11596_ _11596_/A _14969_/Q vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ _13338_/A _13335_/B vssd1 vssd1 vccd1 vccd1 _15131_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10547_ _10548_/A _10548_/B _10548_/C _10548_/D vssd1 vssd1 vccd1 vccd1 _10547_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13266_ _13287_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _15108_/D sky130_fd_sc_hd__nor2_1
X_10478_ _11564_/A _10827_/C _10477_/C _10477_/D vssd1 vssd1 vccd1 vccd1 _10478_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15005_ _15268_/CLK _15005_/D vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__dfxtp_1
X_12217_ _06926_/A _12210_/Y _12212_/Y _12214_/Y _12216_/Y vssd1 vssd1 vccd1 vccd1
+ _12218_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_110_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09376__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13197_ _13404_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _15062_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12148_ _14885_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12148_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12079_ hold2433/X _12099_/A2 _12078_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12079_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08887__B1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08351__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08892__B _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15214_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _08310_/A _08310_/B _08310_/C vssd1 vssd1 vccd1 vccd1 _08312_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08103__A2 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09290_ _09290_/A _09290_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_118_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08241_ _08165_/X _08166_/Y _08164_/Y vssd1 vssd1 vccd1 vccd1 _08242_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_25 _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__B1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_36 _14928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__A _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__B _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08172_/X sky130_fd_sc_hd__or2_1
XANTENNA_58 _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_69 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07123_ _13724_/A1 hold2133/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07614__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12634__S _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10943__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07728__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07054_ _13659_/A1 hold1107/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07054_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10496__C_N _10482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12597__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput165 _15177_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[12] sky130_fd_sc_hd__buf_12
Xoutput176 _15187_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[22] sky130_fd_sc_hd__buf_12
Xoutput187 _15168_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[3] sky130_fd_sc_hd__buf_12
Xoutput198 _14181_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[11] sky130_fd_sc_hd__buf_12
X_07956_ _08014_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _07958_/B sky130_fd_sc_hd__or2_1
XFILLER_0_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06907_ _06907_/A vssd1 vssd1 vccd1 vccd1 _07437_/A sky130_fd_sc_hd__inv_2
X_07887_ _07887_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _07887_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout653_A _15197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08342__A2 _13382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_211_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09557_ _09557_/A _09557_/B _09557_/C vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__and3_2
XANTENNA_fanout820_A _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12809__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11713__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15400_/CLK sky130_fd_sc_hd__clkbuf_16
X_08508_ _08509_/B _08509_/A vssd1 vssd1 vccd1 vccd1 _08508_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10437__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12521__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ _09215_/A _09347_/B _09347_/A vssd1 vssd1 vccd1 vccd1 _09488_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10837__B _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08439_ _09918_/A _13424_/B _13351_/B _08256_/A _08438_/Y vssd1 vssd1 vccd1 vccd1
+ _08440_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _11449_/A _11449_/B _11607_/A _11448_/X vssd1 vssd1 vccd1 vccd1 _11450_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12729__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _10401_/A _10401_/B _10401_/C vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__or3_1
XANTENNA__10275__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11381_ _11381_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13490_/A hold147/X vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__and2_1
XANTENNA__07638__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10332_ _10333_/A _10333_/B _10333_/C vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__and3_2
XFILLER_0_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13051_ _13101_/A _13051_/B vssd1 vssd1 vccd1 vccd1 _13052_/C sky130_fd_sc_hd__or2_1
X_10263_ _10266_/B _10263_/B _10263_/C _10267_/A vssd1 vssd1 vccd1 vccd1 _10265_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11165__A1 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12002_ _12068_/A hold2665/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12002_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11165__B2 _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _10191_/X _10192_/Y _09984_/B _09987_/B vssd1 vssd1 vccd1 vccd1 _10194_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout370 _07899_/Y vssd1 vssd1 vccd1 vccd1 _12260_/A2 sky130_fd_sc_hd__clkbuf_16
Xfanout381 _11943_/S vssd1 vssd1 vccd1 vccd1 _11959_/S sky130_fd_sc_hd__clkbuf_16
Xfanout392 _07879_/X vssd1 vssd1 vccd1 vccd1 _07900_/B sky130_fd_sc_hd__buf_12
XFILLER_0_205_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13953_ _15454_/CLK _13953_/D vssd1 vssd1 vccd1 vccd1 _13953_/Q sky130_fd_sc_hd__dfxtp_1
X_12904_ _13397_/B _13104_/A2 _12903_/X vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _15380_/CLK _13884_/D vssd1 vssd1 vccd1 vccd1 _13884_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12835_ hold921/A _13947_/Q _12915_/S vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12417__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15360_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13404__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ _14348_/Q _14252_/Q _12841_/S vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10979__A1 _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10979__B2 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08192__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14505_ _15440_/CLK _14505_/D vssd1 vssd1 vccd1 vccd1 _14505_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11717_ hold2107/X _13671_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__mux2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11640__A2 _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07844__B2 _15345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ hold937/A hold669/A _14636_/Q _14732_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11648_ _13750_/A _13373_/B _13373_/C _13468_/B _13749_/A vssd1 vssd1 vccd1 vccd1
+ _11648_/X sky130_fd_sc_hd__o32a_1
X_14436_ _15309_/CLK _14436_/D vssd1 vssd1 vccd1 vccd1 _14436_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput12 dmemresp_rdata[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput23 dmemresp_rdata[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 imemresp_data[10] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput45 imemresp_data[20] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
XFILLER_0_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11579_ _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11581_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14367_ _15432_/CLK _14367_/D vssd1 vssd1 vccd1 vccd1 _14367_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10763__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput56 imemresp_data[30] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 in0[11] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_1
Xhold807 hold807/A vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput78 in0[21] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_1
Xinput89 in0[31] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__buf_1
X_13318_ input146/X fanout5/X fanout3/X input114/X vssd1 vssd1 vccd1 vccd1 _13318_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11578__B _14971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold818 hold818/A vssd1 vssd1 vccd1 vccd1 hold818/X sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ _14557_/CLK hold530/X vssd1 vssd1 vccd1 vccd1 hold529/A sky130_fd_sc_hd__dfxtp_1
Xhold829 hold829/A vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08233__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ input151/X fanout6/X fanout4/X input119/X vssd1 vssd1 vccd1 vccd1 _13249_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2208 _07128_/X vssd1 vssd1 vccd1 vccd1 _13938_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2219 _14720_/Q vssd1 vssd1 vccd1 vccd1 hold2219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11594__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ hold885/X _13748_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold886/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2416_A _13749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08790_ _09816_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1507 _13988_/Q vssd1 vssd1 vccd1 vccd1 hold1507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1518 _07615_/X vssd1 vssd1 vccd1 vccd1 _14238_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _15395_/Q vssd1 vssd1 vccd1 vccd1 hold1529/X sky130_fd_sc_hd__dlygate4sd3_1
X_07741_ hold657/X _13714_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold658/A sky130_fd_sc_hd__mux2_1
XANTENNA__12656__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15216__D _15216_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10667__B1 _10666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__B2 _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ hold1861/X _13711_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 _07672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09411_ _09411_/A _09411_/B _09411_/C vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__10762__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12506__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2785_A _11641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15426_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13314__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _11287_/S _09341_/X _09339_/X vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13081__A1 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09273_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09273_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07835__A1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08224_ _08144_/A _08144_/C _08144_/B vssd1 vssd1 vccd1 vccd1 _08226_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08155_ _10873_/A _08702_/B _08209_/A _08155_/D vssd1 vssd1 vccd1 vccd1 _08209_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_16_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout401_A _07477_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07599__A0 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12592__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ _13742_/A1 hold2279/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07106_/X sky130_fd_sc_hd__mux2_1
X_08086_ _08085_/A _08085_/B _08085_/C vssd1 vssd1 vccd1 vccd1 _08088_/D sky130_fd_sc_hd__a21o_1
XANTENNA__08260__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07037_ hold1339/X _13741_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 _07037_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout770_A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13045__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2720 _14838_/Q vssd1 vssd1 vccd1 vccd1 hold2720/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11708__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2731 _15124_/Q vssd1 vssd1 vccd1 vccd1 hold2731/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2742 _15065_/Q vssd1 vssd1 vccd1 vccd1 hold2742/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2753 _15176_/Q vssd1 vssd1 vccd1 vccd1 hold2753/X sky130_fd_sc_hd__dlygate4sd3_1
X_08988_ _14668_/Q _13941_/Q hold881/A _13909_/Q _10425_/S0 _10425_/S1 vssd1 vssd1
+ vccd1 vccd1 _08989_/B sky130_fd_sc_hd__mux4_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07193__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2764 _15063_/Q vssd1 vssd1 vccd1 vccd1 hold2764/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2775 _13020_/X vssd1 vssd1 vccd1 vccd1 _13027_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07939_ hold423/A _14205_/Q hold359/A _14459_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07940_/B sky130_fd_sc_hd__mux4_1
Xhold2786 _15195_/Q vssd1 vssd1 vccd1 vccd1 hold2786/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12112__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2797 _10566_/Y vssd1 vssd1 vccd1 vccd1 _13399_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11009__A _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10950_ _13745_/A1 _12260_/A2 _11514_/B1 _13200_/B _10948_/Y vssd1 vssd1 vccd1 vccd1
+ _10950_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _09606_/Y _09607_/X _09464_/Y _09466_/X vssd1 vssd1 vccd1 vccd1 _09609_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_168_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10881_ _11517_/A _11586_/B _10881_/C _10881_/D vssd1 vssd1 vccd1 vccd1 _10881_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _12620_/A _12620_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__or3b_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07222__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09371__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ _12601_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12552_/C sky130_fd_sc_hd__or2_1
XFILLER_0_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08037__B _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _11507_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/Y sky130_fd_sc_hd__nor2_1
X_12482_ _12482_/A _12482_/B vssd1 vssd1 vccd1 vccd1 _14947_/D sky130_fd_sc_hd__nor2_1
X_15270_ _15270_/CLK _15270_/D vssd1 vssd1 vccd1 vccd1 _15270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11433_ _11575_/A _11434_/C _11434_/A vssd1 vssd1 vccd1 vccd1 _11445_/A sky130_fd_sc_hd__a21oi_1
X_14221_ _15449_/CLK hold104/X vssd1 vssd1 vccd1 vccd1 _14221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10583__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14152_ _15436_/CLK hold702/X vssd1 vssd1 vccd1 vccd1 hold701/A sky130_fd_sc_hd__dfxtp_1
X_11364_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _11563_/A _14956_/Q _14957_/Q _11594_/A vssd1 vssd1 vccd1 vccd1 _10316_/D
+ sky130_fd_sc_hd__a22o_1
X_13103_ _13715_/A1 _13103_/A2 _12330_/X _13203_/B vssd1 vssd1 vccd1 vccd1 _13103_/X
+ sky130_fd_sc_hd__a22o_1
X_14083_ _14083_/CLK _14083_/D vssd1 vssd1 vccd1 vccd1 _14083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11295_ _13594_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__and2_1
XANTENNA__07892__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ hold829/A _13923_/Q _13041_/S vssd1 vssd1 vccd1 vccd1 _13034_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08003__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10246_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10246_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12886__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _10177_/A _10177_/B vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12099__C1 _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12638__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14985_ _15243_/CLK hold148/X vssd1 vssd1 vccd1 vccd1 _14985_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__09503__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12733__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13936_ _14775_/CLK _13936_/D vssd1 vssd1 vccd1 vccd1 _13936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13867_ _14754_/CLK _13867_/D vssd1 vssd1 vccd1 vccd1 _13867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13599__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ _06942_/A _12815_/X _12817_/X vssd1 vssd1 vccd1 vccd1 _12818_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13063__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12497__S0 _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__A _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__B _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _15296_/CLK _13798_/D vssd1 vssd1 vccd1 vccd1 _13798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09362__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12749_ _13879_/Q hold291/A _13847_/Q _13815_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux4_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__B1 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14419_ _14419_/CLK hold548/X vssd1 vssd1 vccd1 vccd1 hold547/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11377__A1 _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ _15436_/CLK hold712/X vssd1 vssd1 vccd1 vccd1 hold711/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__B2 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold604 hold604/A vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 hold615/A vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold626 hold626/A vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold637 hold637/A vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10643__D _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap356 _11460_/B vssd1 vssd1 vccd1 vccd1 _11267_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold648 hold648/A vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09960_ _10166_/A _10338_/B _11536_/B _10166_/C vssd1 vssd1 vccd1 vccd1 _10170_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold659 hold659/A vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08911_ _08794_/A _08794_/B _08794_/C vssd1 vssd1 vccd1 vccd1 _08912_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09891_ _09888_/Y _09889_/X _09734_/B _09734_/Y vssd1 vssd1 vccd1 vccd1 _09892_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12421__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _13929_/Q vssd1 vssd1 vccd1 vccd1 hold2005/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 _13674_/X vssd1 vssd1 vccd1 vccd1 _15381_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 _15270_/Q vssd1 vssd1 vccd1 vccd1 hold2027/X sky130_fd_sc_hd__dlygate4sd3_1
X_08842_ _09117_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _08842_/X sky130_fd_sc_hd__xor2_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2038 _07183_/X vssd1 vssd1 vccd1 vccd1 _13990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12972__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1304 _11839_/X vssd1 vssd1 vccd1 vccd1 _14662_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2049 _13864_/Q vssd1 vssd1 vccd1 vccd1 hold2049/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 _13811_/Q vssd1 vssd1 vccd1 vccd1 hold1315/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__A _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1326 _07781_/X vssd1 vssd1 vccd1 vccd1 _14396_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ hold2691/X _12260_/A2 _12259_/A1 _13185_/B _08771_/Y vssd1 vssd1 vccd1 vccd1
+ _08773_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12629__A1 _13386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1337 _13889_/Q vssd1 vssd1 vccd1 vccd1 hold1337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1348 _07725_/X vssd1 vssd1 vccd1 vccd1 _14344_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 _14364_/Q vssd1 vssd1 vccd1 vccd1 hold1359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13743__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07724_ hold989/X _13730_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold990/A sky130_fd_sc_hd__mux2_1
XANTENNA__12724__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07741__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07655_ hold821/X _13727_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold822/A sky130_fd_sc_hd__mux2_1
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout449_A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _13725_/A1 hold495/X _07593_/S vssd1 vssd1 vccd1 vccd1 hold496/A sky130_fd_sc_hd__mux2_1
XANTENNA__13054__A1 _11287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ _09464_/A _09324_/C _09324_/A vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07808__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _09571_/A _09712_/B _09255_/C _09255_/D vssd1 vssd1 vccd1 vccd1 _09256_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07977__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10__f_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08207_ hold2759/X input30/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13179_/B sky130_fd_sc_hd__mux2_1
X_09187_ _09186_/B _09186_/C _09186_/A vssd1 vssd1 vccd1 vccd1 _09187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07188__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _08901_/A _08893_/A _08926_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08214_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08069_ _08054_/Y _08059_/Y _08068_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08070_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_113_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10100_ _11504_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10100_/Y sky130_fd_sc_hd__nor2_1
X_11080_ _11080_/A _11080_/B vssd1 vssd1 vccd1 vccd1 _11081_/B sky130_fd_sc_hd__or2_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12868__A1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _09852_/A _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _10036_/A sky130_fd_sc_hd__a21bo_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2550 _14829_/Q vssd1 vssd1 vccd1 vccd1 hold2550/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2561 _13579_/X vssd1 vssd1 vccd1 vccd1 _15315_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2572 _13581_/X vssd1 vssd1 vccd1 vccd1 _15316_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2583 _15137_/Q vssd1 vssd1 vccd1 vccd1 hold2583/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2594 _12171_/X vssd1 vssd1 vccd1 vccd1 _14896_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13653__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1860 _07060_/X vssd1 vssd1 vccd1 vccd1 _13876_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1871 _14318_/Q vssd1 vssd1 vccd1 vccd1 hold1871/X sky130_fd_sc_hd__dlygate4sd3_1
X_14770_ _15411_/CLK _14770_/D vssd1 vssd1 vccd1 vccd1 _14770_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ hold1085/X _13671_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__mux2_1
Xhold1882 _11933_/X vssd1 vssd1 vccd1 vccd1 _14753_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1893 _13886_/Q vssd1 vssd1 vccd1 vccd1 hold1893/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07651__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ hold811/X _13721_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 hold812/A sky130_fd_sc_hd__mux2_1
XFILLER_0_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ _15386_/Q hold963/A hold411/A _14390_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _10933_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09151__B _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10864_ _10863_/A _10863_/B _10863_/C vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__a21o_1
X_13652_ hold883/X _13652_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold884/A sky130_fd_sc_hd__mux2_1
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10297__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ hold2732/X _12329_/B _12953_/B1 _13183_/B vssd1 vssd1 vccd1 vccd1 _12603_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10795_/A _10795_/B vssd1 vssd1 vccd1 vccd1 _10814_/A sky130_fd_sc_hd__nand2_1
X_13583_ _10228_/B _13797_/A2 _13582_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _13583_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11901__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10803__B1 _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15324_/CLK _15322_/D vssd1 vssd1 vccd1 vccd1 _15322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12534_ hold1269/X hold2063/X _12560_/S vssd1 vssd1 vccd1 vccd1 _12534_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13401__B _13401_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15253_ _15258_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold153/A sky130_fd_sc_hd__dfxtp_1
X_12465_ hold1735/X hold1531/X _12466_/S vssd1 vssd1 vccd1 vccd1 _12465_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12556__B1 _13149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ _15392_/CLK _14204_/D vssd1 vssd1 vccd1 vccd1 _14204_/Q sky130_fd_sc_hd__dfxtp_1
X_11416_ _11416_/A _11608_/B _11416_/C vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__nand3_1
X_12396_ _15361_/Q _15264_/Q hold935/A _14365_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12396_/X sky130_fd_sc_hd__mux4_1
X_15184_ _15184_/CLK _15184_/D vssd1 vssd1 vccd1 vccd1 _15184_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11347_ _11200_/A _11199_/B _11197_/X vssd1 vssd1 vccd1 vccd1 _11358_/A sky130_fd_sc_hd__a21o_1
X_14135_ _14909_/CLK _14135_/D vssd1 vssd1 vccd1 vccd1 _14135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11278_ _11278_/A _11278_/B _11278_/C vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__nor3_1
X_14066_ _15351_/CLK _14066_/D vssd1 vssd1 vccd1 vccd1 _14066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13017_ _13092_/A1 _13016_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10229_ _10744_/A _09927_/B _09933_/A vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_158_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11531__A1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14968_ _14972_/CLK _14968_/D vssd1 vssd1 vccd1 vccd1 _14968_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12087__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13919_ _15415_/CLK _13919_/D vssd1 vssd1 vccd1 vccd1 _13919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14899_ _14987_/CLK _14899_/D vssd1 vssd1 vccd1 vccd1 _14899_/Q sky130_fd_sc_hd__dfxtp_1
X_07440_ _13240_/A _12607_/A vssd1 vssd1 vccd1 vccd1 _14070_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13036__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ _15346_/Q _14059_/Q vssd1 vssd1 vccd1 vccd1 _07371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10000__B _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ hold405/A _14541_/Q hold987/A _14765_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09110_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11811__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08463__A1 _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ _09979_/B _09864_/A _10022_/A _10183_/A vssd1 vssd1 vccd1 vccd1 _09043_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10270__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10270__B2 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2748_A _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12208__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10654__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold401 hold401/A vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 hold412/A vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold423 hold423/A vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13738__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold434 hold434/A vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 hold445/A vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10951__A _10951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold456 hold456/A vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 hold467/A vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07736__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold478 hold478/A vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 hold489/A vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09943_ _11509_/A _09943_/B vssd1 vssd1 vccd1 vccd1 _09943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout399_A _07577_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _10110_/A _10010_/B _09702_/D _09701_/X vssd1 vssd1 vccd1 vccd1 _09879_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08140__B _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _13992_/Q vssd1 vssd1 vccd1 vccd1 hold1101/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 _11980_/X vssd1 vssd1 vccd1 vccd1 _14799_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08825_ _08825_/A _08825_/B _08825_/C vssd1 vssd1 vccd1 vccd1 _08825_/Y sky130_fd_sc_hd__nand3_2
Xhold1123 _14612_/Q vssd1 vssd1 vccd1 vccd1 hold1123/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _13730_/X vssd1 vssd1 vccd1 vccd1 _15440_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout566_A _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 _15290_/Q vssd1 vssd1 vccd1 vccd1 hold1145/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 _13654_/X vssd1 vssd1 vccd1 vccd1 _15361_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 _14754_/Q vssd1 vssd1 vccd1 vccd1 hold1167/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__B1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ hold459/A _15274_/Q hold927/A _14375_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08756_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08567__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1178 _07177_/X vssd1 vssd1 vccd1 vccd1 _13985_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _14600_/Q vssd1 vssd1 vccd1 vccd1 hold1189/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10089__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07707_ hold531/X _13680_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold532/A sky130_fd_sc_hd__mux2_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _08686_/B _08686_/C _08686_/A vssd1 vssd1 vccd1 vccd1 _08689_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout733_A _14957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07638_ hold903/X _13744_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold904/A sky130_fd_sc_hd__mux2_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11006__B _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07569_ _13396_/A hold161/X vssd1 vssd1 vccd1 vccd1 hold162/A sky130_fd_sc_hd__and2_1
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__A1 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12786__B1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09308_ _09307_/B _09307_/C _09307_/A vssd1 vssd1 vccd1 vccd1 _09308_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10580_ _11507_/A _10577_/X _10579_/X vssd1 vssd1 vccd1 vccd1 _10580_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09239_ _15407_/Q hold693/A _14702_/Q _14766_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09239_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__A _14999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9__f_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12250_ _06926_/A _12243_/Y _12245_/Y _12247_/Y _12249_/Y vssd1 vssd1 vccd1 vccd1
+ _12250_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_181_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12633__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10283__D _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12181_ _12114_/A _12195_/A2 _12180_/X _13491_/A vssd1 vssd1 vccd1 vccd1 _12181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07646__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ hold877/A _13955_/Q hold829/A _13923_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11133_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09427__A _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold990 hold990/A vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _11063_/A _11063_/B _11242_/B vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09801__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2380 _13557_/X vssd1 vssd1 vccd1 vccd1 _15304_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _14840_/CLK _14822_/D vssd1 vssd1 vccd1 vccd1 _14822_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2391 hold2843/X vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__buf_1
XFILLER_0_204_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1690 _06984_/X vssd1 vssd1 vccd1 vccd1 _13803_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08368__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _15394_/CLK _14753_/D vssd1 vssd1 vccd1 vccd1 _14753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ hold1103/X _13654_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11965_/X sky130_fd_sc_hd__mux2_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ hold1719/X _13704_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13704_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _07296_/B _10602_/X _10951_/A vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13018__A1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14684_ _15458_/CLK hold470/X vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11896_ _13651_/A1 hold1603/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_128_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08643__A2_N _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13635_ hold2600/X _13797_/A2 _13634_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15345_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13569__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _10848_/A _10848_/B _10848_/C vssd1 vssd1 vccd1 vccd1 _10847_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11124__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13566_ _14439_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__or2_1
XANTENNA__12872__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10778_ _13711_/A1 _11514_/A2 _11514_/B1 _13199_/B _10776_/Y vssd1 vssd1 vccd1 vccd1
+ _10778_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07410__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15305_ _15305_/CLK _15305_/D vssd1 vssd1 vccd1 vccd1 _15305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12517_ _12692_/A1 _12516_/X _14490_/Q vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08996__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13497_ _13499_/A hold109/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__and2_1
XANTENNA__10474__C _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ _15251_/CLK _15236_/D vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12448_ hold263/A _14303_/Q _14594_/Q _13963_/Q _12460_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12448_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12624__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08748__A2 _13430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15167_ _15365_/CLK _15167_/D vssd1 vssd1 vccd1 vccd1 _15167_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10771__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ _12379_/A _12379_/B _13376_/B vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14118_ _14731_/CLK _14118_/D vssd1 vssd1 vccd1 vccd1 _14118_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11586__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15098_ _15387_/CLK hold754/X vssd1 vssd1 vccd1 vccd1 hold753/A sky130_fd_sc_hd__dfxtp_1
X_06940_ _06940_/A vssd1 vssd1 vccd1 vccd1 _06940_/Y sky130_fd_sc_hd__inv_2
X_14049_ _14105_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08056__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10307__A2 _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10938__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07184__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11806__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08610_ _08610_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _08612_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09590_ _09591_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ _08541_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _08541_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08472_ _08472_/A _08472_/B vssd1 vssd1 vccd1 vccd1 _08511_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07304__B _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08684__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08684__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _07423_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _07423_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09800__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07354_ _07427_/A _07426_/A _07362_/B _07353_/C vssd1 vssd1 vccd1 vccd1 _07904_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_190_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07285_ _08892_/A _08312_/A vssd1 vssd1 vccd1 vccd1 _12254_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09024_ _09661_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09027_/A sky130_fd_sc_hd__and2_1
XANTENNA__11991__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08739__A2 _13386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__B _07974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__S _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 _13693_/A1 vssd1 vssd1 vccd1 vccd1 _13512_/A0 sky130_fd_sc_hd__clkbuf_4
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _15041_/Q vssd1 vssd1 vccd1 vccd1 _13721_/A1 sky130_fd_sc_hd__buf_4
Xfanout722 _14963_/Q vssd1 vssd1 vccd1 vccd1 _11563_/B sky130_fd_sc_hd__buf_6
XFILLER_0_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _14445_/Q _13586_/B _09918_/Y hold2478/X _13579_/C1 vssd1 vssd1 vccd1 vccd1
+ _09926_/X sky130_fd_sc_hd__o221a_1
Xfanout733 _14957_/Q vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__clkbuf_8
Xfanout744 _10304_/C vssd1 vssd1 vccd1 vccd1 _09864_/C sky130_fd_sc_hd__buf_4
Xfanout755 _14950_/Q vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__10929__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 _09542_/A vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__buf_6
XANTENNA__09795__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09857_ _09858_/B _09858_/C _09709_/B _09858_/A vssd1 vssd1 vccd1 vccd1 _09857_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout777 _14944_/Q vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__buf_4
XANTENNA_fanout850_A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 _10351_/A vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__clkbuf_8
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout799 _14490_/Q vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__buf_8
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11716__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _08809_/B _09437_/A _08809_/D _09571_/A vssd1 vssd1 vccd1 vccd1 _08810_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12401__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ _10426_/A _09787_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _09788_/X sky130_fd_sc_hd__o21a_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_104 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ _07900_/B _13386_/B _08669_/X vssd1 vssd1 vccd1 vccd1 _13430_/B sky130_fd_sc_hd__a21oi_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12120__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_115 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__A _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_148 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A1 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ _13703_/A1 hold1633/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__mux2_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__B2 _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10700_/A _11614_/B _10878_/A _10700_/D vssd1 vssd1 vccd1 vccd1 _10702_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11681_ _13745_/A1 hold999/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11681_/X sky130_fd_sc_hd__mux2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13420_ _13440_/S _13420_/B vssd1 vssd1 vccd1 vccd1 _13420_/Y sky130_fd_sc_hd__nand2_1
X_10632_ _10631_/B _10631_/C _10631_/A vssd1 vssd1 vccd1 vccd1 _10633_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_193_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10563_ _10736_/B _10563_/B vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13351_ _13360_/A _13351_/B vssd1 vssd1 vccd1 vccd1 _15142_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _07437_/A _14031_/Q _06935_/Y _15347_/Q vssd1 vssd1 vccd1 vccd1 _12302_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13282_ input133/X fanout6/X fanout4/X input101/X vssd1 vssd1 vccd1 vccd1 _13282_/X
+ sky130_fd_sc_hd__a22o_1
X_10494_ _10494_/A _10494_/B _10494_/C vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__and3_1
XFILLER_0_133_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11687__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15021_ _15188_/CLK _15021_/D vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12233_ _12233_/A _12233_/B vssd1 vssd1 vccd1 vccd1 _12233_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10591__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12931__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12164_ _14893_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__or2_1
XANTENNA__08061__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11115_ _15161_/Q _07812_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _11115_/Y sky130_fd_sc_hd__a21oi_1
X_12095_ hold2418/X _12099_/A2 _12094_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12095_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11046_ _11229_/B _11045_/B _11045_/C vssd1 vssd1 vccd1 vccd1 _11047_/B sky130_fd_sc_hd__a21oi_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09786__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08902__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _15382_/CLK _14805_/D vssd1 vssd1 vccd1 vccd1 _14805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ hold563/X hold849/X hold481/X hold1105/X _12991_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12997_/X sky130_fd_sc_hd__mux4_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14736_ _15444_/CLK _14736_/D vssd1 vssd1 vccd1 vccd1 _14736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11948_ _13703_/A1 hold2267/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09042__D _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08666__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08761__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14667_ _15441_/CLK hold792/X vssd1 vssd1 vccd1 vccd1 hold791/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13098__S0 _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ hold987/X _13700_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold988/A sky130_fd_sc_hd__mux2_1
XANTENNA__13142__A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13618_ _07432_/A _13792_/A2 _13617_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15336_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10485__B _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14598_ _15391_/CLK _14598_/D vssd1 vssd1 vccd1 vccd1 _14598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__A1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ _08179_/B _08441_/B _13548_/X _13178_/A vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _13675_/A1 hold1893/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07070_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15219_ _15222_/CLK _15219_/D vssd1 vssd1 vccd1 vccd1 _15219_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11597__A _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput303 _14846_/Q vssd1 vssd1 vccd1 vccd1 out1[1] sky130_fd_sc_hd__buf_12
XFILLER_0_112_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold2446_A _15459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput314 _14847_/Q vssd1 vssd1 vccd1 vccd1 out1[2] sky130_fd_sc_hd__buf_12
XANTENNA__08277__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput325 _14823_/Q vssd1 vssd1 vccd1 vccd1 out2[10] sky130_fd_sc_hd__buf_12
Xoutput336 _14833_/Q vssd1 vssd1 vccd1 vccd1 out2[20] sky130_fd_sc_hd__buf_12
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput347 _14843_/Q vssd1 vssd1 vccd1 vccd1 out2[30] sky130_fd_sc_hd__buf_12
XFILLER_0_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15219__D _15219_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07972_ _06904_/A _07432_/A _08036_/S vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13022__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _09711_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__and2_2
X_06923_ _06923_/A vssd1 vssd1 vccd1 vccd1 _07453_/A sky130_fd_sc_hd__inv_2
XFILLER_0_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08354__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13317__A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ hold407/A hold533/A hold643/A hold941/A _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09643_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09573_ _09864_/A _09712_/B _09573_/C _09573_/D vssd1 vssd1 vccd1 vccd1 _09573_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12438__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08521_/X _08524_/B _08524_/C vssd1 vssd1 vccd1 vccd1 _08571_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12453__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ hold319/A hold831/A hold959/A hold561/A _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08456_/B sky130_fd_sc_hd__mux4_1
XANTENNA__08752__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12367__S _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout431_A _11763_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout529_A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13052__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07406_ hold262/X _13317_/A vssd1 vssd1 vccd1 vccd1 _14036_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08386_ _09661_/A _09437_/A vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__and2_1
XFILLER_0_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07880__A2 _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07337_ _07903_/C _09344_/B _07336_/Y vssd1 vssd1 vccd1 vccd1 _07337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10826__D _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _08569_/A vssd1 vssd1 vccd1 vccd1 _07328_/B sky130_fd_sc_hd__inv_2
XFILLER_0_147_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09007_ _09136_/A _09714_/C _09864_/D _09009_/A vssd1 vssd1 vccd1 vccd1 _09011_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07199_ hold1443/X _13519_/A0 _07214_/S vssd1 vssd1 vccd1 vccd1 _07199_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A2 _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout530 _08869_/A vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__clkbuf_8
Xfanout541 _08763_/S1 vssd1 vssd1 vccd1 vccd1 _08868_/S1 sky130_fd_sc_hd__clkbuf_8
X_09909_ _10071_/A _10071_/B vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__nor2_1
Xfanout552 _11316_/S1 vssd1 vssd1 vccd1 vccd1 _11306_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout563 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _12198_/S sky130_fd_sc_hd__clkbuf_4
Xfanout574 _11501_/S0 vssd1 vssd1 vccd1 vccd1 _11506_/S0 sky130_fd_sc_hd__buf_8
XANTENNA__12141__A1 hold2628/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 _10166_/C vssd1 vssd1 vccd1 vccd1 _11542_/B sky130_fd_sc_hd__clkbuf_8
Xfanout596 _09979_/C vssd1 vssd1 vccd1 vccd1 _10827_/D sky130_fd_sc_hd__clkbuf_4
X_12920_ _12920_/A _12920_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07225__A _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12951_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12852_/C sky130_fd_sc_hd__or2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13661__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11802_ hold1493/X _13656_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 _11802_/X sky130_fd_sc_hd__mux2_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13641__A1 _08253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12782_ _13171_/A _12782_/B vssd1 vssd1 vccd1 vccd1 _14959_/D sky130_fd_sc_hd__nor2_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11101__C1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _15421_/CLK hold350/X vssd1 vssd1 vccd1 vccd1 hold349/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09940__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11733_ hold479/X hold2813/X _11745_/S vssd1 vssd1 vccd1 vccd1 hold480/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07879__B _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _15426_/CLK _14452_/D vssd1 vssd1 vccd1 vccd1 _14452_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ _13728_/A1 hold2259/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _13404_/A _13403_/B vssd1 vssd1 vccd1 vccd1 _15194_/D sky130_fd_sc_hd__and2_1
X_10615_ _10461_/A _10461_/B _10454_/Y vssd1 vssd1 vccd1 vccd1 _10631_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14383_ _15090_/CLK _14383_/D vssd1 vssd1 vccd1 vccd1 _14383_/Q sky130_fd_sc_hd__dfxtp_1
X_11595_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11601_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__A0 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ input88/X fanout2/X _13333_/X vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ _10543_/Y _10544_/X _10370_/Y _10373_/X vssd1 vssd1 vccd1 vccd1 _10548_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output183_A _15194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13265_ input94/X fanout1/X _13264_/X vssd1 vssd1 vccd1 vccd1 _13266_/B sky130_fd_sc_hd__a21oi_1
X_10477_ _11564_/A _10827_/C _10477_/C _10477_/D vssd1 vssd1 vccd1 vccd1 _10477_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_122_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15004_ _15004_/CLK hold708/X vssd1 vssd1 vccd1 vccd1 _15004_/Q sky130_fd_sc_hd__dfxtp_1
X_12216_ _12243_/A _12215_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _12216_/Y sky130_fd_sc_hd__o21ai_1
X_13196_ _13397_/A _13196_/B vssd1 vssd1 vccd1 vccd1 _15061_/D sky130_fd_sc_hd__and2_1
XANTENNA__08584__B1 _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12380__A1 _13174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12740__S _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ hold2634/X _12173_/A2 _12146_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_209_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12078_ _14979_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12078_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11029_ _10814_/B _10817_/B _11027_/Y _11028_/X vssd1 vssd1 vccd1 vccd1 _11029_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__10143__B1 _14957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12976__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14719_ _15045_/CLK _14719_/D vssd1 vssd1 vccd1 vccd1 _14719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08243_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_15 _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_26 _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__A1 _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_37 _14935_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08244_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_48 _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__B _12288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12915__S _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_59 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07122_ _13690_/A1 hold1711/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07122_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07075__A0 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08811__A1 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07053_ _13691_/A1 hold1889/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07053_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13699__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07378__A1 _15342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput166 _15178_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[13] sky130_fd_sc_hd__buf_12
XFILLER_0_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput177 _15188_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[23] sky130_fd_sc_hd__buf_12
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13746__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput188 _15169_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[4] sky130_fd_sc_hd__buf_12
Xoutput199 _14182_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_wdata[12] sky130_fd_sc_hd__buf_12
XFILLER_0_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07955_ _08312_/A _08075_/B _07952_/Y _08010_/A vssd1 vssd1 vccd1 vccd1 _07956_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout381_A _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout479_A _06959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ _13241_/A vssd1 vssd1 vccd1 vccd1 _07438_/A sky130_fd_sc_hd__inv_2
X_07886_ _12254_/A _12254_/B _07889_/C vssd1 vssd1 vccd1 vccd1 _07887_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__or2_1
XFILLER_0_210_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout646_A _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _09555_/B _09555_/C _09555_/A vssd1 vssd1 vccd1 vccd1 _09557_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_210_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08507_ _08507_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _08509_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout813_A _14489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _09775_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09491_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_210_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10837__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ hold2670/X _11643_/B _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08438_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08369_ _08877_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _08369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ _11288_/A1 _13398_/B _10259_/X vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__a21o_2
X_11380_ _11564_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _11381_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08604__A _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10328_/X _10329_/Y _10151_/X _10156_/B vssd1 vssd1 vccd1 vccd1 _10333_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12126__A _15003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ _10600_/B _10601_/A vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__or2_1
X_13050_ _13046_/X _13047_/X _13049_/X _13048_/X _13050_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _13051_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11165__A2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _12063_/A _12001_/B vssd1 vssd1 vccd1 vccd1 _14813_/D sky130_fd_sc_hd__and2_1
XANTENNA__13656__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__C _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10193_ _09984_/B _09987_/B _10191_/X _10192_/Y vssd1 vssd1 vccd1 vccd1 _10193_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__12560__S _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07654__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout360 _12326_/Y vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__buf_12
XFILLER_0_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout371 _12252_/B vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__buf_8
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout382 _11960_/S vssd1 vssd1 vccd1 vccd1 _11943_/S sky130_fd_sc_hd__clkbuf_16
Xfanout393 _07745_/Y vssd1 vssd1 vccd1 vccd1 _07761_/S sky130_fd_sc_hd__clkbuf_16
X_13952_ _15453_/CLK _13952_/D vssd1 vssd1 vccd1 vccd1 _13952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ _13674_/A1 _13103_/A2 _13078_/B1 _13195_/B vssd1 vssd1 vccd1 vccd1 _12903_/X
+ sky130_fd_sc_hd__a22o_1
X_13883_ _15379_/CLK _13883_/D vssd1 vssd1 vccd1 vccd1 _13883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11904__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _15448_/Q _13915_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12834_/X sky130_fd_sc_hd__mux2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ hold583/X _14124_/Q _12841_/S vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__mux2_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10979__A2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14504_ _15268_/CLK _14504_/D vssd1 vssd1 vccd1 vccd1 _14504_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11716_ hold549/X _13736_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 hold550/A sky130_fd_sc_hd__mux2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ hold845/A hold947/A _15084_/Q _14377_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12696_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_72_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14435_ _15305_/CLK _14435_/D vssd1 vssd1 vccd1 vccd1 _14435_/Q sky130_fd_sc_hd__dfxtp_1
X_11647_ _11479_/A _11483_/X _11644_/Y _11645_/X vssd1 vssd1 vccd1 vccd1 _13373_/C
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__12735__S _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 dmemresp_rdata[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12050__A0 hold2555/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput24 dmemresp_rdata[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput35 imemresp_data[11] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
X_14366_ _15265_/CLK _14366_/D vssd1 vssd1 vccd1 vccd1 _14366_/Q sky130_fd_sc_hd__dfxtp_1
Xinput46 imemresp_data[21] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
X_11578_ _11578_/A _14971_/Q _11578_/C vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__and3_1
Xinput57 imemresp_data[31] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput68 in0[12] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _13317_/A _13317_/B vssd1 vssd1 vccd1 vccd1 _15125_/D sky130_fd_sc_hd__nor2_1
Xhold808 hold808/A vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 in0[22] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10529_ _11517_/A _11564_/B _10696_/A _10528_/D vssd1 vssd1 vccd1 vccd1 _10530_/C
+ sky130_fd_sc_hd__a22o_1
Xhold819 hold819/A vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14297_ _15456_/CLK _14297_/D vssd1 vssd1 vccd1 vccd1 _14297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08233__B _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13248_ _13287_/A _13248_/B vssd1 vssd1 vccd1 vccd1 _15102_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _13386_/A _13179_/B vssd1 vssd1 vccd1 vccd1 _15044_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08652__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2209 _13899_/Q vssd1 vssd1 vccd1 vccd1 hold2209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11594__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1508 _07180_/X vssd1 vssd1 vccd1 vccd1 _13988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1519 _15370_/Q vssd1 vssd1 vccd1 vccd1 hold1519/X sky130_fd_sc_hd__dlygate4sd3_1
X_07740_ hold629/X _13746_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold630/A sky130_fd_sc_hd__mux2_1
XFILLER_0_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10116__B1 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12656__A2 _13153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07671_ hold1837/X hold2764/X _07676_/S vssd1 vssd1 vccd1 vccd1 _07671_/X sky130_fd_sc_hd__mux2_1
X_09410_ _09411_/A _09411_/B _09411_/C vssd1 vssd1 vccd1 vccd1 _09410_/X sky130_fd_sc_hd__and3_1
XFILLER_0_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11814__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10762__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09341_ _09341_/A _09341_/B vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__xor2_1
XANTENNA_hold2778_A _09342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12813__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15232__D _15232_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_89_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _09274_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_132_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08223_ _08222_/B _08222_/C _08222_/A vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07739__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08154_ _10873_/A _08702_/B _08209_/A _08155_/D vssd1 vssd1 vccd1 vccd1 _08156_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12592__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _13741_/A1 hold2117/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07105_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08085_ _08085_/A _08085_/B _08085_/C vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_147_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07036_ hold685/X _13674_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold686/A sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout596_A _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2710 _15165_/Q vssd1 vssd1 vccd1 vccd1 hold2710/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2721 _12050_/X vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2732 _15048_/Q vssd1 vssd1 vccd1 vccd1 hold2732/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _08989_/A _08987_/B vssd1 vssd1 vccd1 vccd1 _08987_/Y sky130_fd_sc_hd__nor2_1
Xhold2743 _15177_/Q vssd1 vssd1 vccd1 vccd1 hold2743/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2754 _15120_/Q vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2765 hold2765/A vssd1 vssd1 vccd1 vccd1 hold2765/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ _08197_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07938_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10107__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2776 _13027_/X vssd1 vssd1 vccd1 vccd1 hold2776/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2787 _15102_/Q vssd1 vssd1 vccd1 vccd1 hold2787/X sky130_fd_sc_hd__buf_1
XFILLER_0_199_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2798 _14216_/Q vssd1 vssd1 vccd1 vccd1 hold2798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11009__B _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ _14085_/Q _07867_/X _11996_/C _07865_/X vssd1 vssd1 vccd1 vccd1 _07869_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11724__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _09464_/Y _09466_/X _09606_/Y _09607_/X vssd1 vssd1 vccd1 vccd1 _09608_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09702__B _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ _11351_/B _11564_/B _11614_/B _11541_/A vssd1 vssd1 vccd1 vccd1 _10881_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__nand2_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07222__B _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ _12546_/X _12547_/X _12549_/X _12548_/X _06943_/Y _12700_/S1 vssd1 vssd1
+ vccd1 vccd1 _12551_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_176_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09371__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ hold227/A _14329_/Q hold557/A _13989_/Q _11501_/S0 _11501_/S1 vssd1 vssd1
+ vccd1 vccd1 _11502_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ _08179_/A _08637_/B _13146_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12482_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12032__A0 hold2471/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ _15445_/CLK _14220_/D vssd1 vssd1 vccd1 vccd1 _14220_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07649__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _11431_/A _11574_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11434_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _15438_/CLK _14151_/D vssd1 vssd1 vccd1 vccd1 _14151_/Q sky130_fd_sc_hd__dfxtp_1
X_11363_ _11524_/B _11361_/X _11254_/B _11254_/Y vssd1 vssd1 vccd1 vccd1 _11364_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _13102_/A _13102_/B _13102_/C vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__and3_1
X_10314_ _11594_/A _11563_/A _14956_/Q _14957_/Q vssd1 vssd1 vccd1 vccd1 _10483_/A
+ sky130_fd_sc_hd__nand4_2
X_14082_ _15425_/CLK _14082_/D vssd1 vssd1 vccd1 vccd1 _14082_/Q sky130_fd_sc_hd__dfxtp_1
X_11294_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _13371_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08539__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13532__A0 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ _15419_/Q _14554_/Q hold513/A _14778_/Q _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13033_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07892__B _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10245_ _10426_/A _10242_/X _10244_/X _10255_/A1 vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12219__B_N _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _09816_/A _10338_/D _09968_/A _09965_/X vssd1 vssd1 vccd1 vccd1 _10177_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14984_ _14987_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 _14984_/Q sky130_fd_sc_hd__dfxtp_4
X_13935_ _15436_/CLK _13935_/D vssd1 vssd1 vccd1 vccd1 _13935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13866_ _15394_/CLK _13866_/D vssd1 vssd1 vccd1 vccd1 _13866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ _12917_/A1 _12816_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09267__A1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13797_ hold2600/X _13797_/A2 _13634_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15426_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08228__B _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__S1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09362__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ hold223/A hold637/A _14606_/Q _13975_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12748_/X sky130_fd_sc_hd__mux4_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10821__A1 _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__B2 _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12465__S _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ _13388_/B _12325_/B _12678_/X vssd1 vssd1 vccd1 vccd1 _12679_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_167_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13150__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14418_ _15093_/CLK hold898/X vssd1 vssd1 vccd1 vccd1 hold897/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15398_ _15398_/CLK _15398_/D vssd1 vssd1 vccd1 vccd1 _15398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11377__A2 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14349_ _14612_/CLK _14349_/D vssd1 vssd1 vccd1 vccd1 _14349_/Q sky130_fd_sc_hd__dfxtp_1
Xhold605 hold605/A vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold616 hold616/A vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 hold627/A vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold649 hold649/A vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08910_ _08909_/B _08909_/C _08909_/A vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11809__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2526_A _15354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ _09734_/B _09734_/Y _09888_/Y _09889_/X vssd1 vssd1 vccd1 vccd1 _09995_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_111_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 _07119_/X vssd1 vssd1 vccd1 vccd1 _13929_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12421__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08841_ _08841_/A _08841_/B vssd1 vssd1 vccd1 vccd1 _08842_/B sky130_fd_sc_hd__nand2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 _14719_/Q vssd1 vssd1 vccd1 vccd1 hold2017/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2028 _13512_/X vssd1 vssd1 vccd1 vccd1 _15270_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 _14273_/Q vssd1 vssd1 vccd1 vccd1 hold2039/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 _13810_/Q vssd1 vssd1 vccd1 vccd1 hold1305/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _06992_/X vssd1 vssd1 vccd1 vccd1 _13811_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1327 _15383_/Q vssd1 vssd1 vccd1 vccd1 hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__B _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ hold2726/X input5/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13185_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12629__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1338 _07073_/X vssd1 vssd1 vccd1 vccd1 _13889_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 _13890_/Q vssd1 vssd1 vccd1 vccd1 hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07723_ hold1109/X _13729_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 _07723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07654_ hold1161/X _13693_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 _07654_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07585_ _15044_/Q hold801/X _07593_/S vssd1 vssd1 vccd1 vccd1 hold802/A sky130_fd_sc_hd__mux2_1
XANTENNA__13054__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08138__B _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _09324_/A _09464_/A _09324_/C vssd1 vssd1 vccd1 vccd1 _09324_/X sky130_fd_sc_hd__or3_1
XFILLER_0_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09255_ _09571_/A _09866_/B _09255_/C _09255_/D vssd1 vssd1 vccd1 vccd1 _09255_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout511_A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout609_A _15208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__A0 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ _12252_/B _08206_/B vssd1 vssd1 vccd1 vccd1 _08206_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ _09186_/A _09186_/B _09186_/C vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08137_ _08893_/A _08926_/A _08809_/B _08901_/A vssd1 vssd1 vccd1 vccd1 _08139_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08864__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07993__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08564_/A1 _08061_/Y _08063_/Y _08065_/Y _08067_/Y vssd1 vssd1 vccd1 vccd1
+ _08068_/X sky130_fd_sc_hd__o32a_1
XANTENNA_fanout880_A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11719__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07019_ hold1029/X _13657_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07019_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10030_ _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10038_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10423__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2540 _15356_/Q vssd1 vssd1 vccd1 vccd1 _08535_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2551 _12032_/X vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2562 _14987_/Q vssd1 vssd1 vccd1 vccd1 hold2562/X sky130_fd_sc_hd__buf_2
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2573 _15317_/Q vssd1 vssd1 vccd1 vccd1 _10228_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2584 _08045_/X vssd1 vssd1 vccd1 vccd1 _08046_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2595 _15346_/Q vssd1 vssd1 vccd1 vccd1 _13241_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1850 _07081_/X vssd1 vssd1 vccd1 vccd1 _13894_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1861 _14293_/Q vssd1 vssd1 vccd1 vccd1 hold1861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1872 _07698_/X vssd1 vssd1 vccd1 vccd1 _14318_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11981_ hold455/X _13736_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 hold456/A sky130_fd_sc_hd__mux2_1
Xhold1883 _14325_/Q vssd1 vssd1 vccd1 vccd1 hold1883/X sky130_fd_sc_hd__dlygate4sd3_1
X_13720_ hold1669/X hold2376/X _13732_/S vssd1 vssd1 vccd1 vccd1 _13720_/X sky130_fd_sc_hd__mux2_1
Xhold1894 _07070_/X vssd1 vssd1 vccd1 vccd1 _13886_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10932_ _11493_/A _10929_/X _10931_/X vssd1 vssd1 vccd1 vccd1 _10932_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ hold917/X _13651_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold918/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09249__A1 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _10863_/A _10863_/B _10863_/C vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10297__C _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12602_ _13027_/A _12602_/B _12602_/C vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__and3_1
XFILLER_0_137_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13582_ _14447_/Q _13634_/B vssd1 vssd1 vccd1 vccd1 _13582_/X sky130_fd_sc_hd__or2_1
XFILLER_0_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10817_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15321_ _15325_/CLK _15321_/D vssd1 vssd1 vccd1 vccd1 _15321_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10803__A1 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12533_ hold711/X hold749/X hold579/X hold1521/X _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12533_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10803__B2 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15252_ _15258_/CLK hold134/X vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__dfxtp_1
X_12464_ hold1559/X hold2802/X _14144_/Q hold2241/X _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12464_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ _14750_/CLK hold498/X vssd1 vssd1 vccd1 vccd1 hold497/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12556__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13753__B1 _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11415_ _11174_/A _11174_/C _11174_/B vssd1 vssd1 vccd1 vccd1 _11416_/C sky130_fd_sc_hd__a21bo_1
X_15183_ _15190_/CLK _15183_/D vssd1 vssd1 vccd1 vccd1 _15183_/Q sky130_fd_sc_hd__dfxtp_2
X_12395_ _12395_/A _12395_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__or3b_1
XANTENNA__08999__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14134_ _14485_/CLK _14134_/D vssd1 vssd1 vccd1 vccd1 _14134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11346_ _11346_/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14065_ _15351_/CLK _14065_/D vssd1 vssd1 vccd1 vccd1 _14065_/Q sky130_fd_sc_hd__dfxtp_1
X_11277_ _11278_/A _11278_/B _11278_/C vssd1 vssd1 vccd1 vccd1 _11280_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ hold1095/X hold667/X _13041_/S vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10414__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _10744_/A _10228_/B vssd1 vssd1 vccd1 vccd1 _10401_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08003__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11531__A2 _15227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10159_ _10156_/X _10157_/Y _10041_/X _10046_/B vssd1 vssd1 vccd1 vccd1 _10160_/C
+ sky130_fd_sc_hd__a211o_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14967_ _14971_/CLK _14967_/D vssd1 vssd1 vccd1 vccd1 _14967_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10769__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13145__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ _15451_/CLK _13918_/D vssd1 vssd1 vccd1 vccd1 _13918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14898_ _15250_/CLK _14898_/D vssd1 vssd1 vccd1 vccd1 _14898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13849_ _15439_/CLK hold566/X vssd1 vssd1 vccd1 vccd1 hold565/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07370_ _15346_/Q _14059_/Q vssd1 vssd1 vccd1 vccd1 _07370_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09660__A1 _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09040_ _09571_/A _09860_/A _08887_/X _08888_/X _09858_/A vssd1 vssd1 vccd1 vccd1
+ _09045_/A sky130_fd_sc_hd__a32o_1
XANTENNA__10270__A2 _14964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09099__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10654__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold402 hold402/A vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold413/A vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 hold424/A vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 hold435/A vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08702__A _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 hold446/A vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold457 hold457/A vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold468 hold468/A vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _09514_/A _09939_/X _09941_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _09943_/B
+ sky130_fd_sc_hd__o211a_1
Xhold479 hold479/A vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__buf_1
XFILLER_0_102_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09873_ _10115_/A _10115_/B _09724_/C _09724_/D _09727_/B vssd1 vssd1 vccd1 vccd1
+ _09881_/A sky130_fd_sc_hd__a41o_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07726__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08825_/A _08825_/B _08825_/C vssd1 vssd1 vccd1 vccd1 _08824_/X sky130_fd_sc_hd__and3_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _07185_/X vssd1 vssd1 vccd1 vccd1 _13992_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 _14111_/Q vssd1 vssd1 vccd1 vccd1 hold1113/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _11787_/X vssd1 vssd1 vccd1 vccd1 _14612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 _14014_/Q vssd1 vssd1 vccd1 vccd1 hold1135/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07752__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1146 _13532_/X vssd1 vssd1 vccd1 vccd1 _15290_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1157 _14471_/Q vssd1 vssd1 vccd1 vccd1 hold1157/X sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _08981_/A _08752_/X _08754_/X vssd1 vssd1 vccd1 vccd1 _08755_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout461_A _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 _11934_/X vssd1 vssd1 vccd1 vccd1 _14754_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1179 _14751_/Q vssd1 vssd1 vccd1 vccd1 hold1179/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ hold317/X _13679_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold318/A sky130_fd_sc_hd__mux2_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _08686_/A _08686_/B _08686_/C vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__nand3_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ hold433/X _13743_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold434/A sky130_fd_sc_hd__mux2_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout726_A _14960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11006__C _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _13396_/A hold155/X vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__and2_1
XFILLER_0_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09307_ _09307_/A _09307_/B _09307_/C vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__and3_2
XANTENNA__11589__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07499_ hold1863/X _13738_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07499_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09651__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07199__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ _09514_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _09238_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__A1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09169_ _09979_/B _09712_/A _10022_/B _10183_/A vssd1 vssd1 vccd1 vccd1 _09171_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12633__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11200_ _11200_/A _11200_/B vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09708__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _14901_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _11504_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11131_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12134__A _14878_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold980 hold980/A vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold991 hold991/A vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07228__A _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _11517_/A _11620_/B _11062_/C _11242_/A vssd1 vssd1 vccd1 vccd1 _11242_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13664__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _10013_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__xor2_2
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07662__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2370 hold2853/X vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__buf_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14821_ _14840_/CLK _14821_/D vssd1 vssd1 vccd1 vccd1 _14821_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2381 _15328_/Q vssd1 vssd1 vccd1 vccd1 _07345_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2392 _13553_/X vssd1 vssd1 vccd1 vccd1 _15302_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10589__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1680 _07518_/X vssd1 vssd1 vccd1 vccd1 _14143_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _15397_/CLK _14752_/D vssd1 vssd1 vccd1 vccd1 _14752_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1691 _14307_/Q vssd1 vssd1 vccd1 vccd1 hold1691/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11964_ hold1945/X _13653_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08059__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ hold879/X _13703_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold880/A sky130_fd_sc_hd__mux2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ hold2751/X _10914_/Y _11283_/S vssd1 vssd1 vccd1 vccd1 _10915_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14683_ _15068_/CLK hold488/X vssd1 vssd1 vccd1 vccd1 hold487/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11895_ _11928_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__or2_4
XFILLER_0_169_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11912__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13634_ input43/X _13634_/B vssd1 vssd1 vccd1 vccd1 _13634_/X sky130_fd_sc_hd__or2_1
X_10846_ _10660_/A _10660_/C _10660_/B vssd1 vssd1 vccd1 vccd1 _10848_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__13423__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12321__S0 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11124__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _08966_/A _09222_/B _13564_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _13565_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13412__B _13412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777_ hold2772/X input20/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12872__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ _15304_/CLK _15304_/D vssd1 vssd1 vccd1 vccd1 _15304_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07410__B _07410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12516_ hold461/A hold733/A _12560_/S vssd1 vssd1 vccd1 vccd1 _12516_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13496_ _13499_/A hold99/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__and2_1
XFILLER_0_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12529__A1 _13382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10474__D _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _15243_/CLK _15235_/D vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12447_ _14786_/Q hold789/A _14626_/Q _14722_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12447_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12624__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15166_ _15365_/CLK _15166_/D vssd1 vssd1 vccd1 vccd1 _15166_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12378_ _12377_/X _12364_/X _12601_/A vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _15438_/CLK _14117_/D vssd1 vssd1 vccd1 vccd1 _14117_/Q sky130_fd_sc_hd__dfxtp_1
X_11329_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__or2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15097_ _15289_/CLK hold412/X vssd1 vssd1 vccd1 vccd1 hold411/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14048_ _14105_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08056__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10938__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08668__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A1 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08381__B2 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08540_ _09918_/A _12270_/B _13352_/B _08256_/A _08539_/Y vssd1 vssd1 vccd1 vccd1
+ _08541_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08133__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2593_A _14992_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ _09858_/B _08383_/B _08470_/X vssd1 vssd1 vccd1 vccd1 _08472_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_175_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08684__A2 _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11822__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _07422_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12768__A1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2760_A _15191_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12312__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07353_ hold2655/X _07362_/B _07353_/C _07353_/D vssd1 vssd1 vccd1 vccd1 _07910_/B
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__B1 _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15240__D _15240_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11440__A1 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07284_ _08892_/A _08312_/A vssd1 vssd1 vccd1 vccd1 _07889_/C sky130_fd_sc_hd__and2_1
XFILLER_0_31_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09023_ _09816_/A _09676_/D vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07747__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout701 _15046_/Q vssd1 vssd1 vccd1 vccd1 _13693_/A1 sky130_fd_sc_hd__buf_4
Xfanout712 _13687_/A1 vssd1 vssd1 vccd1 vccd1 _13654_/A1 sky130_fd_sc_hd__clkbuf_4
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ hold2477/X _09925_/A2 _13590_/B _09922_/Y _09924_/X vssd1 vssd1 vccd1 vccd1
+ _09925_/X sky130_fd_sc_hd__a2111o_1
Xfanout723 _14962_/Q vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__clkbuf_8
Xfanout734 _11537_/A vssd1 vssd1 vccd1 vccd1 _09724_/C sky130_fd_sc_hd__buf_4
XANTENNA__12153__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _10304_/C vssd1 vssd1 vccd1 vccd1 _09714_/C sky130_fd_sc_hd__clkbuf_4
Xfanout756 _14950_/Q vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10929__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _09856_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__xnor2_1
Xfanout767 _14947_/Q vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__buf_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout778 _08908_/A vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__buf_4
XANTENNA__09795__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 _14941_/Q vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__clkbuf_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07482__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__A1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ _08674_/A _08673_/A _08673_/B vssd1 vssd1 vccd1 vccd1 _08812_/A sky130_fd_sc_hd__o21bai_2
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _13883_/Q hold621/A hold397/A _13819_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09787_/X sky130_fd_sc_hd__mux4_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ _13671_/A1 hold2031/X _07010_/S vssd1 vssd1 vccd1 vccd1 _06999_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_198_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ hold2451/X _08526_/B _08846_/C _08737_/Y _08735_/X vssd1 vssd1 vccd1 vccd1
+ _13386_/B sky130_fd_sc_hd__a221o_4
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12456__B1 _13145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_105 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_127 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_149 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _13663_/A1 _12260_/A2 _12259_/A1 _13184_/B _08667_/Y vssd1 vssd1 vccd1 vccd1
+ _08669_/X sky130_fd_sc_hd__a221o_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11732__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _10700_/A _11614_/B _10878_/A _10700_/D vssd1 vssd1 vccd1 vccd1 _10878_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _13711_/A1 hold1513/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11680_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _10631_/A _10631_/B _10631_/C vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_165_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10234__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ _13360_/A _13350_/B vssd1 vssd1 vccd1 vccd1 _15141_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ _10562_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10563_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_146_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _12301_/A _12301_/B _12301_/C _12308_/A vssd1 vssd1 vccd1 vccd1 _12326_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13659__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _13287_/A _13281_/B vssd1 vssd1 vccd1 vccd1 _15113_/D sky130_fd_sc_hd__nor2_1
X_10493_ _10320_/A _10320_/C _10320_/B vssd1 vssd1 vccd1 vccd1 _10494_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15020_ _15184_/CLK _15020_/D vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07657__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _13863_/Q _13991_/Q _12237_/S vssd1 vssd1 vccd1 vccd1 _12233_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12931__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ hold2509/X _12173_/A2 _12162_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12163_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11114_ _13590_/A _11113_/C _11113_/A vssd1 vssd1 vccd1 vccd1 _11114_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_208_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _14987_/Q _12096_/B _12096_/C _12124_/D vssd1 vssd1 vccd1 vccd1 _12094_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__09235__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11907__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ _11229_/B _11045_/B _11045_/C vssd1 vssd1 vccd1 vccd1 _11047_/A sky130_fd_sc_hd__and3_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09786__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _15408_/CLK _14804_/D vssd1 vssd1 vccd1 vccd1 _14804_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ hold1365/X hold1609/X hold553/X hold1967/X _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12996_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _15087_/CLK _14735_/D vssd1 vssd1 vccd1 vccd1 _14735_/Q sky130_fd_sc_hd__dfxtp_1
X_11947_ _13735_/A1 hold863/X _11959_/S vssd1 vssd1 vccd1 vccd1 hold864/A sky130_fd_sc_hd__mux2_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _15405_/CLK hold598/X vssd1 vssd1 vccd1 vccd1 hold597/A sky130_fd_sc_hd__dfxtp_1
X_11878_ hold737/X _15052_/Q _11893_/S vssd1 vssd1 vccd1 vccd1 hold738/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13098__S1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13617_ input34/X _13636_/B vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__or2_1
XFILLER_0_157_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10829_ _11564_/A _11537_/B _10830_/C _10830_/D vssd1 vssd1 vccd1 vccd1 _10829_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__10258__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14597_ _15435_/CLK _14597_/D vssd1 vssd1 vccd1 vccd1 _14597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10485__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13548_ _14430_/Q _13554_/B vssd1 vssd1 vccd1 vccd1 _13548_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13479_ _13479_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _15238_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15218_ _15222_/CLK _15218_/D vssd1 vssd1 vccd1 vccd1 _15218_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09379__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__B _14968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput304 _14865_/Q vssd1 vssd1 vccd1 vccd1 out1[20] sky130_fd_sc_hd__buf_12
XANTENNA__08252__A _08253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput315 _14875_/Q vssd1 vssd1 vccd1 vccd1 out1[30] sky130_fd_sc_hd__buf_12
XANTENNA__08277__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput326 _14824_/Q vssd1 vssd1 vccd1 vccd1 out2[11] sky130_fd_sc_hd__buf_12
XFILLER_0_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput337 _14834_/Q vssd1 vssd1 vccd1 vccd1 out2[21] sky130_fd_sc_hd__buf_12
XFILLER_0_168_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _15313_/CLK _15149_/D vssd1 vssd1 vccd1 vccd1 _15149_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput348 _14844_/Q vssd1 vssd1 vccd1 vccd1 out2[31] sky130_fd_sc_hd__buf_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold2439_A _14990_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _07921_/A _07920_/A _07920_/B vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__13022__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ _10129_/A _09709_/B _09709_/C _09709_/D vssd1 vssd1 vccd1 vccd1 _09711_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11817__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06922_ _06922_/A vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__inv_2
XANTENNA__12686__B1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _10246_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_207_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12221__B _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15235__D _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09572_ _09864_/A _09712_/B _09573_/C _09573_/D vssd1 vssd1 vccd1 vccd1 _09572_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__10022__A _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08523_ _08524_/C _08524_/B vssd1 vssd1 vccd1 vccd1 _08523_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12533__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _12241_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13089__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07405_ _07405_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14035_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_190_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08385_ _08312_/A _09437_/A _08312_/D _08309_/X vssd1 vssd1 vccd1 vccd1 _08397_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A _11961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11413__A1 _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _07812_/A _07812_/B vssd1 vssd1 vccd1 vccd1 _07336_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07267_ _10024_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__and2_1
XANTENNA__10692__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ _09006_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_130_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07198_ hold713/X _13666_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold714/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12913__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13469__A2 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _15426_/Q vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__buf_6
XANTENNA__11727__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 _08869_/A vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__clkbuf_8
Xfanout542 _15423_/Q vssd1 vssd1 vccd1 vccd1 _08763_/S1 sky130_fd_sc_hd__buf_8
X_09908_ _09905_/X _09906_/Y _09751_/X _09754_/X vssd1 vssd1 vccd1 vccd1 _10071_/B
+ sky130_fd_sc_hd__a211oi_2
Xfanout553 _15423_/Q vssd1 vssd1 vccd1 vccd1 _11316_/S1 sky130_fd_sc_hd__buf_4
Xfanout564 _07822_/S vssd1 vssd1 vccd1 vccd1 _07816_/S sky130_fd_sc_hd__buf_8
Xfanout575 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _11501_/S0 sky130_fd_sc_hd__clkbuf_8
Xfanout586 _15216_/Q vssd1 vssd1 vccd1 vccd1 _10166_/C sky130_fd_sc_hd__buf_4
X_09839_ _09839_/A _09839_/B _09839_/C vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__or3_1
Xfanout597 _15212_/Q vssd1 vssd1 vccd1 vccd1 _09979_/C sky130_fd_sc_hd__buf_6
XANTENNA__12772__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07225__B _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _12846_/X _12847_/X _12849_/X _12848_/X _12950_/S0 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12851_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_198_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ hold521/X _13655_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold522/A sky130_fd_sc_hd__mux2_1
XANTENNA__12524__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _13106_/A1 _13158_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12782_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_185_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09845__A1 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09845__B2 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14926_/CLK hold850/X vssd1 vssd1 vccd1 vccd1 hold849/A sky130_fd_sc_hd__dfxtp_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _13718_/A1 hold1989/X _11745_/S vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__mux2_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__A _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09940__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07241__A _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _15320_/CLK _14451_/D vssd1 vssd1 vccd1 vccd1 _14451_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_193_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11663_ _13727_/A1 hold1223/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11663_/X sky130_fd_sc_hd__mux2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13402_ _13479_/A _13402_/B vssd1 vssd1 vccd1 vccd1 _15193_/D sky130_fd_sc_hd__and2_1
XFILLER_0_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10614_ _10614_/A _10614_/B vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__xnor2_1
X_14382_ _15089_/CLK _14382_/D vssd1 vssd1 vccd1 vccd1 _14382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ _11594_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ input152/X fanout6/A fanout4/A input120/X vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10545_ _10370_/Y _10373_/X _10543_/Y _10544_/X vssd1 vssd1 vccd1 vccd1 _10548_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_88_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_130_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15445_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ input158/X fanout6/X fanout4/X input126/X vssd1 vssd1 vccd1 vccd1 _13264_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10476_ _11564_/A _10827_/C _10477_/C _10477_/D vssd1 vssd1 vccd1 vccd1 _10476_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15003_ _15258_/CLK hold172/X vssd1 vssd1 vccd1 vccd1 _15003_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output176_A _15187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12904__A1 _13397_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12215_ _15390_/Q hold439/A _14685_/Q _14749_/Q _12198_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12215_/X sky130_fd_sc_hd__mux4_1
X_13195_ _13397_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _15060_/D sky130_fd_sc_hd__and2_1
XFILLER_0_209_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08584__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08584__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__A2 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _14884_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13418__A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ hold2495/X _12099_/A2 _12076_/X _13492_/A vssd1 vssd1 vccd1 vccd1 _12077_/X
+ sky130_fd_sc_hd__o211a_1
X_11028_ _11027_/A _11027_/B _11014_/Y vssd1 vssd1 vccd1 vccd1 _11028_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10143__A1 _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10143__B2 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12979_ _10741_/X _13104_/A2 _12978_/X vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__a21o_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13153__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14718_ _15428_/CLK _14718_/D vssd1 vssd1 vccd1 vccd1 _14718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14649_ _15421_/CLK hold364/X vssd1 vssd1 vccd1 vccd1 hold363/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_16 _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_27 _14921_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08170_ _08102_/A _07323_/C _08029_/X _08169_/X _08496_/A vssd1 vssd1 vccd1 vccd1
+ _08172_/B sky130_fd_sc_hd__a311o_1
XANTENNA_38 _14935_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _15235_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07121_ _13689_/A1 hold1805/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07121_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15278_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08811__A2 _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07052_ _13657_/A1 hold1997/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput167 _15179_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[14] sky130_fd_sc_hd__buf_12
XFILLER_0_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput178 _15189_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[24] sky130_fd_sc_hd__buf_12
Xoutput189 _15170_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[5] sky130_fd_sc_hd__buf_12
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ _07952_/Y _08010_/A _08312_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08014_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12123__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06905_ _06905_/A vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__inv_2
XFILLER_0_208_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07885_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _11287_/S sky130_fd_sc_hd__nand2_4
Xclkbuf_leaf_188_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _14595_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07760__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _09555_/A _09555_/B _09555_/C vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__nand3_2
XANTENNA__09827__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12378__S _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10687__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ _08507_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _08616_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ hold2641/X _09344_/B _09346_/B vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__12831__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07933__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10837__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _08437_/A _08437_/B vssd1 vssd1 vccd1 vccd1 _13351_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout806_A _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08368_ _14662_/Q _13935_/Q _15436_/Q _13903_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08369_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_191_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ _08340_/A _08378_/A _10951_/A _07319_/D vssd1 vssd1 vccd1 vccd1 _07321_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_112_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15448_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08604__B _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ _10151_/X _10156_/B _10328_/X _10329_/Y vssd1 vssd1 vccd1 vccd1 _10333_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12126__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07000__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10261_ _10600_/B _10601_/A vssd1 vssd1 vccd1 vccd1 _10261_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12841__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ _12066_/A hold2676/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10192_ _10191_/B _10191_/C _10191_/A vssd1 vssd1 vccd1 vccd1 _10192_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08661__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__A _15357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout361 _07390_/A vssd1 vssd1 vccd1 vccd1 _09494_/A1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07236__A _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 _10433_/A vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_179_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _14754_/CLK sky130_fd_sc_hd__clkbuf_16
X_13951_ _14419_/CLK _13951_/D vssd1 vssd1 vccd1 vccd1 _13951_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout383 _11895_/X vssd1 vssd1 vccd1 vccd1 _11911_/S sky130_fd_sc_hd__buf_12
XFILLER_0_199_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11322__B1 _07900_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout394 _07745_/Y vssd1 vssd1 vccd1 vccd1 _07777_/S sky130_fd_sc_hd__buf_12
XANTENNA__13672__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _13102_/A _12902_/B _12902_/C vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__and3_1
X_13882_ _15089_/CLK _13882_/D vssd1 vssd1 vccd1 vccd1 _13882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07670__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ hold1813/X _14546_/Q hold2811/X hold1439/X _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12833_/X sky130_fd_sc_hd__mux4_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09170__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12764_ hold673/X _14220_/Q hold305/A hold587/A _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12764_/X sky130_fd_sc_hd__mux4_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11715_ hold1447/X _13669_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14503_ _14791_/CLK _14503_/D vssd1 vssd1 vccd1 vccd1 _14503_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ _12695_/A _12695_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__or3b_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11920__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ _11644_/Y _11645_/X _11479_/A _11483_/X vssd1 vssd1 vccd1 vccd1 _13373_/B
+ sky130_fd_sc_hd__o211a_1
X_14434_ _15305_/CLK _14434_/D vssd1 vssd1 vccd1 vccd1 _14434_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 dmemresp_rdata[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14365_ _15072_/CLK _14365_/D vssd1 vssd1 vccd1 vccd1 _14365_/Q sky130_fd_sc_hd__dfxtp_1
Xinput25 dmemresp_rdata[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13420__B _13420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput36 imemresp_data[12] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11577_ _11577_/A _14970_/Q vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_103_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _15382_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 imemresp_data[22] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_109_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13316_ input81/X fanout2/X _13315_/X vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput58 imemresp_data[3] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput69 in0[13] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
X_10528_ _11517_/A _11564_/B _10696_/A _10528_/D vssd1 vssd1 vccd1 vccd1 _10696_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold809 hold809/A vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ _15287_/CLK _14296_/D vssd1 vssd1 vccd1 vccd1 _14296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13247_ input76/X fanout1/X _13246_/X vssd1 vssd1 vccd1 vccd1 _13248_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08006__B1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10459_ _11594_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _10460_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13178_ _13178_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _15043_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08652__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12129_ hold2523/X _12129_/A2 _12128_/X _12063_/A vssd1 vssd1 vccd1 vccd1 _12129_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13148__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1509 _15278_/Q vssd1 vssd1 vccd1 vccd1 hold1509/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12105__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10116__B2 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07670_ hold1311/X _11921_/A0 _07676_/S vssd1 vssd1 vccd1 vccd1 _07670_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07580__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12198__S _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09340_ _09340_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09341_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10300__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10001__A2_N _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ _09271_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11830__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ _08222_/A _08222_/B _08222_/C vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08153_ _08152_/A _08152_/B _08152_/C vssd1 vssd1 vccd1 vccd1 _08155_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12227__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11131__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ _13740_/A1 hold1743/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07104_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08084_ _08312_/A _08012_/B _08012_/D _08009_/X vssd1 vssd1 vccd1 vccd1 _08085_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07035_ hold1277/X _13673_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 _07035_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07755__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12975__S0 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10355__B2 _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2700 _14834_/Q vssd1 vssd1 vccd1 vccd1 hold2700/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout589_A _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2711 _15184_/Q vssd1 vssd1 vccd1 vccd1 hold2711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2722 _14841_/Q vssd1 vssd1 vccd1 vccd1 hold2722/X sky130_fd_sc_hd__dlygate4sd3_1
X_08986_ hold757/A _14217_/Q hold605/A _14471_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08987_/B sky130_fd_sc_hd__mux4_1
Xhold2733 _08568_/X vssd1 vssd1 vccd1 vccd1 hold2733/X sky130_fd_sc_hd__buf_1
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2744 _15179_/Q vssd1 vssd1 vccd1 vccd1 hold2744/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2755 _15168_/Q vssd1 vssd1 vccd1 vccd1 hold2755/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ hold595/A _14237_/Q hold381/A _14109_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07938_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2766 _12980_/Y vssd1 vssd1 vccd1 vccd1 _13166_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2777 _15118_/Q vssd1 vssd1 vccd1 vccd1 _09338_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10107__B2 _13195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2788 _15104_/Q vssd1 vssd1 vccd1 vccd1 hold2788/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A _14950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2799 _14759_/Q vssd1 vssd1 vccd1 vccd1 hold2799/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11855__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ _14093_/Q _14092_/Q _14083_/Q vssd1 vssd1 vccd1 vccd1 _11996_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07490__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09607_ _09604_/Y _09605_/X _09421_/Y _09461_/A vssd1 vssd1 vccd1 vccd1 _09607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09702__C _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07799_ hold643/X _13737_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold644/A sky130_fd_sc_hd__mux2_1
XFILLER_0_210_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ _09442_/A _09441_/B _09439_/X vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ _09466_/X _09467_/Y _09323_/Y _09328_/B vssd1 vssd1 vccd1 vccd1 _09471_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11740__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ _11510_/A1 _11493_/Y _11495_/Y _11497_/Y _11499_/Y vssd1 vssd1 vccd1 vccd1
+ _11500_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12480_ _12327_/A _12479_/X _12477_/X vssd1 vssd1 vccd1 vccd1 _13146_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_136_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _11431_/A _11574_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14150_ _14731_/CLK hold556/X vssd1 vssd1 vccd1 vccd1 hold555/A sky130_fd_sc_hd__dfxtp_1
X_11362_ _11254_/B _11254_/Y _11524_/B _11361_/X vssd1 vssd1 vccd1 vccd1 _11364_/A
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__10594__A1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _13101_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _13102_/C sky130_fd_sc_hd__or2_1
X_10313_ _10033_/A _11588_/B _10117_/B _10115_/X vssd1 vssd1 vccd1 vccd1 _10318_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13667__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14081_ _15293_/CLK _14081_/D vssd1 vssd1 vccd1 vccd1 _14081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11293_ _11107_/A _11112_/B _11481_/A vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__a21bo_1
X_13032_ _13107_/A _13032_/B vssd1 vssd1 vccd1 vccd1 _14969_/D sky130_fd_sc_hd__nor2_1
XANTENNA__07665__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _10244_/A _10244_/B vssd1 vssd1 vccd1 vccd1 _10244_/X sky130_fd_sc_hd__or2_1
XANTENNA__07892__C _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__xnor2_1
X_14983_ _15248_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 _14983_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11915__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13934_ _15437_/CLK _13934_/D vssd1 vssd1 vccd1 vccd1 _13934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ _15397_/CLK _13865_/D vssd1 vssd1 vccd1 vccd1 _13865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ hold407/A hold533/A _12841_/S vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13796_ hold2641/X _13797_/A2 _13632_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15425_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12747_ _14798_/Q _14510_/Q hold351/A _14734_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12747_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10821__A2 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12678_ _13665_/A1 _13103_/A2 _13078_/B1 _13186_/B vssd1 vssd1 vccd1 vccd1 _12678_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11629_ _11629_/A _11629_/B vssd1 vssd1 vccd1 vccd1 _11630_/B sky130_fd_sc_hd__xnor2_1
X_14417_ _15196_/CLK hold842/X vssd1 vssd1 vccd1 vccd1 hold841/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13150__B _13150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15397_ _15397_/CLK hold520/X vssd1 vssd1 vccd1 vccd1 hold519/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14348_ _15410_/CLK _14348_/D vssd1 vssd1 vccd1 vccd1 _14348_/Q sky130_fd_sc_hd__dfxtp_1
Xhold606 hold606/A vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold617 hold617/A vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 hold628/A vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14279_ _14602_/CLK _14279_/D vssd1 vssd1 vccd1 vccd1 _14279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold639 hold639/A vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08840_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__nor2_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _14531_/Q vssd1 vssd1 vccd1 vccd1 hold2007/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2018 _11898_/X vssd1 vssd1 vccd1 vccd1 _14719_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _14234_/Q vssd1 vssd1 vccd1 vccd1 hold2029/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _06991_/X vssd1 vssd1 vccd1 vccd1 _13810_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _12252_/B _08771_/B vssd1 vssd1 vccd1 vccd1 _08771_/Y sky130_fd_sc_hd__nor2_1
Xhold1317 _14597_/Q vssd1 vssd1 vccd1 vccd1 hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 _13676_/X vssd1 vssd1 vccd1 vccd1 _15383_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 _13854_/Q vssd1 vssd1 vccd1 vccd1 hold1339/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11825__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07722_ hold631/X _13728_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold632/A sky130_fd_sc_hd__mux2_1
XANTENNA__11298__C1 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07653_ hold379/X _13659_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold380/A sky130_fd_sc_hd__mux2_1
XFILLER_0_177_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07584_ _13690_/A1 hold2093/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07584_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09323_ _09324_/A _09464_/A _09324_/C vssd1 vssd1 vccd1 vccd1 _09323_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08138__C _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13341__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _09571_/A _09866_/B _09255_/C _09255_/D vssd1 vssd1 vccd1 vccd1 _09254_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08435__A _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08205_ _08190_/Y _08195_/Y _08204_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08206_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ _09184_/B _09184_/C _09184_/A vssd1 vssd1 vccd1 vccd1 _09186_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout504_A _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__A1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ _13690_/A1 _12260_/A2 _12259_/A1 _13178_/B _08134_/Y vssd1 vssd1 vccd1 vccd1
+ _08136_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08864__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12391__S _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _08869_/A _08066_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _08067_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ hold1025/X _13656_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12948__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout873_A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10423__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2530 _15032_/Q vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2541 hold2860/X vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2552 _14453_/Q vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__buf_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2563 _12161_/X vssd1 vssd1 vccd1 vccd1 _14891_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08969_ _08969_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__xnor2_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2574 _13583_/X vssd1 vssd1 vccd1 vccd1 _15317_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11735__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1840 _07055_/X vssd1 vssd1 vccd1 vccd1 _13871_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2585 _08047_/X vssd1 vssd1 vccd1 vccd1 _14428_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11828__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1851 _14117_/Q vssd1 vssd1 vccd1 vccd1 hold1851/X sky130_fd_sc_hd__dlygate4sd3_1
X_11980_ hold1111/X _13669_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__mux2_1
Xhold2596 _15162_/Q vssd1 vssd1 vccd1 vccd1 _11297_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1862 _07672_/X vssd1 vssd1 vccd1 vccd1 _14293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1873 _13983_/Q vssd1 vssd1 vccd1 vccd1 hold1873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1884 _07705_/X vssd1 vssd1 vccd1 vccd1 _14325_/D sky130_fd_sc_hd__dlygate4sd3_1
X_10931_ _11504_/A _10930_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _10931_/X sky130_fd_sc_hd__o21a_1
Xhold1895 _14555_/Q vssd1 vssd1 vccd1 vccd1 hold1895/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_116_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _11566_/A _15222_/Q vssd1 vssd1 vccd1 vccd1 _10863_/C sky130_fd_sc_hd__and2_1
X_13650_ _13683_/A _13650_/B vssd1 vssd1 vccd1 vccd1 _13650_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12601_ _12601_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _12602_/C sky130_fd_sc_hd__or2_1
XFILLER_0_184_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12253__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13581_ _09927_/B _13586_/B _13580_/Y _13797_/C1 vssd1 vssd1 vccd1 vccd1 _13581_/X
+ sky130_fd_sc_hd__o211a_1
X_10793_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10793_/X sky130_fd_sc_hd__and2b_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12566__S _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13251__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12607_/A _12532_/B vssd1 vssd1 vccd1 vccd1 _14949_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08552__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15320_ _15320_/CLK _15320_/D vssd1 vssd1 vccd1 vccd1 _15320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10803__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08345__A _08345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ _12642_/B1 _12458_/X _12462_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12470_/A
+ sky130_fd_sc_hd__o211a_1
X_15251_ _15251_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10016__B1 _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ _11569_/A _11605_/B _11414_/C _11608_/A vssd1 vssd1 vccd1 vccd1 _11608_/B
+ sky130_fd_sc_hd__nand4_2
X_14202_ _15390_/CLK _14202_/D vssd1 vssd1 vccd1 vccd1 _14202_/Q sky130_fd_sc_hd__dfxtp_1
X_15182_ _15184_/CLK _15182_/D vssd1 vssd1 vccd1 vccd1 _15182_/Q sky130_fd_sc_hd__dfxtp_2
X_12394_ _12644_/A1 _12389_/X _12393_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12395_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_73_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__B _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ _14776_/CLK hold760/X vssd1 vssd1 vccd1 vccd1 hold759/A sky130_fd_sc_hd__dfxtp_1
X_11345_ _11567_/A _15227_/Q vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14064_ _15351_/CLK _14064_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12939__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ _11468_/B _11276_/B vssd1 vssd1 vccd1 vccd1 _11278_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11516__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output256_A _14430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ hold1079/X hold1625/X _13041_/S vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12713__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10227_ _11288_/A1 _13397_/B _10107_/X vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_88_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10414__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10158_ _10041_/X _10046_/B _10156_/X _10157_/Y vssd1 vssd1 vccd1 vccd1 _10160_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_131_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14966_ _14971_/CLK _14966_/D vssd1 vssd1 vccd1 vccd1 _14966_/Q sky130_fd_sc_hd__dfxtp_4
X_10089_ _09941_/A _10086_/X _10088_/X vssd1 vssd1 vccd1 vccd1 _10089_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_11_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09115__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13145__B _13145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13917_ _15450_/CLK _13917_/D vssd1 vssd1 vccd1 vccd1 _13917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12492__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14897_ _15250_/CLK _14897_/D vssd1 vssd1 vccd1 vccd1 _14897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_146_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13848_ _15087_/CLK hold664/X vssd1 vssd1 vccd1 vccd1 hold663/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08448__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ hold269/X vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10000__D _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09660__A2 _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15449_ _15449_/CLK _15449_/D vssd1 vssd1 vccd1 vccd1 _15449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09099__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11755__A0 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 hold403/A vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 hold414/A vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 hold425/A vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold436 hold436/A vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08702__B _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold447 hold447/A vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold458 hold458/A vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09941_/X sky130_fd_sc_hd__or2_1
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15238__D _15238_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09872_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _09888_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08823_ _08820_/Y _08821_/X _08710_/Y _08714_/B vssd1 vssd1 vccd1 vccd1 _08825_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08923__B2 _14950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _14784_/Q vssd1 vssd1 vccd1 vccd1 hold1103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _07483_/X vssd1 vssd1 vccd1 vccd1 _14111_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _14314_/Q vssd1 vssd1 vccd1 vccd1 hold1125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 _07207_/X vssd1 vssd1 vccd1 vccd1 _14014_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _08989_/A _08753_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08754_/X sky130_fd_sc_hd__o21a_1
Xhold1147 _14021_/Q vssd1 vssd1 vccd1 vccd1 hold1147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 _11668_/X vssd1 vssd1 vccd1 vccd1 _14471_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _14124_/Q vssd1 vssd1 vccd1 vccd1 hold1169/X sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ hold1883/X _13744_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 _07705_/X sky130_fd_sc_hd__mux2_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08685_ _08908_/A _09026_/B _08685_/C _09712_/A vssd1 vssd1 vccd1 vccd1 _08686_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout454_A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _15004_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ hold567/X _11921_/A0 _07642_/S vssd1 vssd1 vccd1 vccd1 hold568/A sky130_fd_sc_hd__mux2_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07567_ _13396_/A hold193/X vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__and2_1
XANTENNA_fanout621_A _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__D _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09305_/B _09305_/C _09305_/A vssd1 vssd1 vccd1 vccd1 _09307_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07498_ hold941/X _13737_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 hold942/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09237_ _14670_/Q _13943_/Q hold723/A _13911_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09238_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13735__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ _09714_/A _10129_/A _09003_/X _09004_/X _10126_/A vssd1 vssd1 vccd1 vccd1
+ _09173_/A sky130_fd_sc_hd__a32o_1
XANTENNA__11746__A0 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08119_ _15364_/Q _15267_/Q _15075_/Q _14368_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08119_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09708__B _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ hold767/A _15277_/Q hold943/A _14378_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09099_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13010__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ hold813/A _14231_/Q hold825/A _14485_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11131_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold970 hold970/A vssd1 vssd1 vccd1 vccd1 hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/A vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _11517_/A _11620_/B _11062_/C _11242_/A vssd1 vssd1 vccd1 vccd1 _11063_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12397__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold992 hold992/A vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _10013_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__nor2_1
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2360 _14996_/Q vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__buf_2
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _14840_/CLK _14820_/D vssd1 vssd1 vccd1 vccd1 _14820_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2371 _13569_/X vssd1 vssd1 vccd1 vccd1 _15310_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2382 hold2834/X vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__buf_1
XFILLER_0_203_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2393 _15031_/Q vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07244__A _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1670 _13720_/X vssd1 vssd1 vccd1 vccd1 _15430_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1681 _13909_/Q vssd1 vssd1 vccd1 vccd1 hold1681/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14751_ _15429_/CLK _14751_/D vssd1 vssd1 vccd1 vccd1 _14751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1692 _07687_/X vssd1 vssd1 vccd1 vccd1 _14307_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11963_ hold1797/X _13652_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 _11963_/X sky130_fd_sc_hd__mux2_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15383_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13680__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ hold1607/X _13735_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13702_/X sky130_fd_sc_hd__mux2_1
X_10914_ _10958_/B _10914_/B vssd1 vssd1 vccd1 vccd1 _10914_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ hold571/X _13715_/A1 _11894_/S vssd1 vssd1 vccd1 vccd1 hold572/A sky130_fd_sc_hd__mux2_1
X_14682_ _15292_/CLK hold878/X vssd1 vssd1 vccd1 vccd1 hold877/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10845_ _10844_/B _10844_/C _10844_/A vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__a21o_1
X_13633_ hold2641/X _13797_/A2 _13632_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15344_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12321__S1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _14438_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13564_/X sky130_fd_sc_hd__or2_1
X_10776_ _11320_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _15305_/CLK _15303_/D vssd1 vssd1 vccd1 vccd1 _15303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12515_ hold409/A _14114_/Q _12560_/S vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13495_ _13495_/A hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__and2_1
XFILLER_0_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ hold893/A _15266_/Q _15074_/Q _14367_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12446_/X sky130_fd_sc_hd__mux4_1
X_15234_ _15243_/CLK _15234_/D vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08803__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08602__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15165_ _15365_/CLK _15165_/D vssd1 vssd1 vccd1 vccd1 _15165_/Q sky130_fd_sc_hd__dfxtp_2
X_12377_ _12700_/S1 _12366_/X _12370_/X _12376_/X vssd1 vssd1 vccd1 vccd1 _12377_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11328_ _11328_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11463_/A sky130_fd_sc_hd__nor2_1
X_14116_ _14955_/CLK hold562/X vssd1 vssd1 vccd1 vccd1 hold561/A sky130_fd_sc_hd__dfxtp_1
X_15096_ _15385_/CLK hold554/X vssd1 vssd1 vccd1 vccd1 hold553/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14047_ _14105_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__dfxtp_1
X_11259_ _11329_/A _11258_/C _11258_/A vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08381__A2 _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13156__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14949_ _15222_/CLK _14949_/D vssd1 vssd1 vccd1 vccd1 _14949_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08669__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15455_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ _08893_/A _09858_/A _09858_/B _08901_/A vssd1 vssd1 vccd1 vccd1 _08470_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ _07812_/A _07903_/C _07450_/B _11650_/B vssd1 vssd1 vccd1 vccd1 _14051_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_159_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12217__A1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09618__C1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07352_ _15340_/Q _15339_/Q _15338_/Q _15332_/Q vssd1 vssd1 vccd1 vccd1 _07353_/C
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12312__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__B2 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07283_ _07283_/A _07283_/B vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11440__A2 _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12934__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _08915_/A _08914_/B _08914_/A vssd1 vssd1 vccd1 vccd1 _09035_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_127_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09809__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__B1 _10259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _14445_/Q _09923_/B _10082_/B _07390_/A vssd1 vssd1 vccd1 vccd1 _09924_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout702 _13659_/A1 vssd1 vssd1 vccd1 vccd1 _13725_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout713 hold2376/X vssd1 vssd1 vccd1 vccd1 _13687_/A1 sky130_fd_sc_hd__buf_4
Xfanout724 _14962_/Q vssd1 vssd1 vccd1 vccd1 _10108_/C sky130_fd_sc_hd__buf_2
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout735 _14956_/Q vssd1 vssd1 vccd1 vccd1 _11537_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07763__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout746 _14953_/Q vssd1 vssd1 vccd1 vccd1 _10304_/C sky130_fd_sc_hd__clkbuf_4
X_09855_ _09856_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__nand2b_1
Xfanout757 _14949_/Q vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__buf_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 _10700_/A vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__clkbuf_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_A _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout779 _14944_/Q vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__buf_6
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout669_A _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _08806_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ hold201/A _14319_/Q _14610_/Q _13979_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09786_/X sky130_fd_sc_hd__mux4_1
X_06998_ _13703_/A1 hold1237/X _07010_/S vssd1 vssd1 vccd1 vccd1 _06998_/X sky130_fd_sc_hd__mux2_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08737_ _07320_/B _10024_/A _08570_/Y _12258_/S vssd1 vssd1 vccd1 vccd1 _08737_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12456__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_106 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14973_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout836_A _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ hold2743/X input4/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__mux2_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07619_ hold733/X _13725_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 hold734/A sky130_fd_sc_hd__mux2_1
XANTENNA__07883__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _08500_/A _08500_/C _08500_/B vssd1 vssd1 vccd1 vccd1 _08610_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10630_ _10795_/B _10629_/C _10629_/A vssd1 vssd1 vccd1 vccd1 _10631_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07003__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10561_ _10559_/X _10561_/B vssd1 vssd1 vccd1 vccd1 _10736_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ _07437_/A _14086_/Q _07875_/X _12299_/X vssd1 vssd1 vccd1 vccd1 _12301_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13708__A1 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13280_ input68/X fanout1/X _13279_/X vssd1 vssd1 vccd1 vccd1 _13281_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10492_ _10491_/B _10491_/C _10491_/A vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ _12231_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_122_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__A1 _11564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12392__B1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__A _15226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12931__A2 _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _14892_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13675__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _11113_/A _13590_/A _11113_/C vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__and3_1
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12093_ hold2420/X _12099_/A2 _12092_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09235__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11044_ _10863_/B _10863_/C _10863_/A vssd1 vssd1 vccd1 vccd1 _11045_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2190 _11830_/X vssd1 vssd1 vccd1 vccd1 _14653_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _15380_/CLK hold794/X vssd1 vssd1 vccd1 vccd1 hold793/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _14077_/CLK sky130_fd_sc_hd__clkbuf_16
X_12995_ _12995_/A _12995_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__or3b_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11923__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14734_ _15278_/CLK _14734_/D vssd1 vssd1 vccd1 vccd1 _14734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _13734_/A1 hold2101/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__mux2_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _15372_/CLK hold998/X vssd1 vssd1 vccd1 vccd1 hold997/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ hold1015/X _13698_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_139_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13616_ _07431_/A _13792_/A2 _13615_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15335_/D
+ sky130_fd_sc_hd__o211a_1
X_10828_ _14954_/Q _10827_/C _10827_/D _14953_/Q vssd1 vssd1 vccd1 vccd1 _10830_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14596_ _15264_/CLK _14596_/D vssd1 vssd1 vccd1 vccd1 _14596_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11958__A0 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10485__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07626__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13547_ hold443/X _08441_/B _13546_/X _13178_/A vssd1 vssd1 vccd1 vccd1 _15299_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10759_ _11504_/A _10758_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _10759_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_124_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13478_ _13487_/A hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__and2_1
XFILLER_0_180_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15217_ _15222_/CLK _15217_/D vssd1 vssd1 vccd1 vccd1 _15217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12429_ _13378_/B _12325_/B _12428_/X vssd1 vssd1 vccd1 vccd1 _12429_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput305 _14866_/Q vssd1 vssd1 vccd1 vccd1 out1[21] sky130_fd_sc_hd__buf_12
XFILLER_0_140_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput316 _14876_/Q vssd1 vssd1 vccd1 vccd1 out1[31] sky130_fd_sc_hd__buf_12
Xoutput327 _14825_/Q vssd1 vssd1 vccd1 vccd1 out2[12] sky130_fd_sc_hd__buf_12
Xoutput338 _14835_/Q vssd1 vssd1 vccd1 vccd1 out2[22] sky130_fd_sc_hd__buf_12
X_15148_ _15309_/CLK _15148_/D vssd1 vssd1 vccd1 vccd1 _15148_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput349 _14816_/Q vssd1 vssd1 vccd1 vccd1 out2[3] sky130_fd_sc_hd__buf_12
XFILLER_0_61_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ _09918_/A _13412_/B vssd1 vssd1 vccd1 vccd1 _07970_/Y sky130_fd_sc_hd__nor2_1
X_15079_ _15079_/CLK _15079_/D vssd1 vssd1 vccd1 vccd1 _15079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07583__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ _06921_/A vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__inv_2
XANTENNA__09364__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12686__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_0_clk/A
+ sky130_fd_sc_hd__clkbuf_16
X_09640_ _10426_/A _09637_/X _09639_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09641_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10303__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09571_ _09571_/A _09714_/A _09714_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _09573_/D
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12438__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10022__B _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _14083_/CLK sky130_fd_sc_hd__clkbuf_16
X_08522_ _08335_/B _08335_/C _08428_/B _08380_/A vssd1 vssd1 vccd1 vccd1 _08524_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10449__B1 _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11833__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12533__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08453_ _12247_/A _08450_/X _08452_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _08454_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07404_ _07404_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14034_/D sky130_fd_sc_hd__nor2_1
X_08384_ _08384_/A _08498_/A vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_190_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07335_ _07903_/C _07359_/A vssd1 vssd1 vccd1 vccd1 _07812_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11413__A2 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout417_A _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07758__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ _11605_/A _10306_/A vssd1 vssd1 vccd1 vccd1 _07267_/B sky130_fd_sc_hd__or2_1
XFILLER_0_6_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10692__B _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ _10126_/A _09004_/X _09003_/X vssd1 vssd1 vccd1 vccd1 _09006_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_116_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07197_ hold1853/X _13665_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12374__B1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout786_A _14941_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout510 _10252_/A vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__buf_4
XANTENNA__07493__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 _08880_/A1 vssd1 vssd1 vccd1 vccd1 _08564_/A1 sky130_fd_sc_hd__clkbuf_8
X_09907_ _09751_/X _09754_/X _09905_/X _09906_/Y vssd1 vssd1 vccd1 vccd1 _10071_/A
+ sky130_fd_sc_hd__o211a_1
Xfanout532 _08869_/A vssd1 vssd1 vccd1 vccd1 _08873_/A sky130_fd_sc_hd__buf_4
Xfanout543 _12211_/S1 vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__clkbuf_8
Xfanout554 _11501_/S1 vssd1 vssd1 vccd1 vccd1 _10930_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout565 _08275_/S0 vssd1 vssd1 vccd1 vccd1 _07822_/S sky130_fd_sc_hd__buf_8
XANTENNA__08976__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 _15422_/Q vssd1 vssd1 vccd1 vccd1 _08275_/S0 sky130_fd_sc_hd__buf_8
X_09838_ _09835_/Y _09836_/X _09684_/Y _09686_/X vssd1 vssd1 vccd1 vccd1 _09839_/C
+ sky130_fd_sc_hd__o211a_1
Xfanout587 _11536_/B vssd1 vssd1 vccd1 vccd1 _11378_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__12772__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout598 _11588_/A vssd1 vssd1 vccd1 vccd1 _10827_/C sky130_fd_sc_hd__buf_4
XFILLER_0_198_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12429__A1 _13378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09769_ _12221_/B _09767_/Y _09914_/C _08526_/B hold2773/X vssd1 vssd1 vccd1 vccd1
+ _09769_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_198_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _14956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11743__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11800_ hold923/X _13654_/A1 _11812_/S vssd1 vssd1 vccd1 vccd1 hold924/A sky130_fd_sc_hd__mux2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12524__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ _13080_/A1 _12779_/X _12777_/X vssd1 vssd1 vccd1 vccd1 _13158_/B sky130_fd_sc_hd__a21oi_4
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09845__A2 _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11731_ _15037_/Q hold439/X _11745_/S vssd1 vssd1 vccd1 vccd1 hold440/A sky130_fd_sc_hd__mux2_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07241__B _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _15320_/CLK _14450_/D vssd1 vssd1 vccd1 vccd1 _14450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _13693_/A1 hold2109/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13401_ _13404_/A _13401_/B vssd1 vssd1 vccd1 vccd1 _15192_/D sky130_fd_sc_hd__and2_1
X_10613_ _10614_/A _10614_/B vssd1 vssd1 vccd1 vccd1 _10794_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11593_ _11445_/B _11593_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14381_ _15056_/CLK _14381_/D vssd1 vssd1 vccd1 vccd1 _14381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07668__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13332_ _13338_/A _13332_/B vssd1 vssd1 vccd1 vccd1 _15130_/D sky130_fd_sc_hd__nor2_1
X_10544_ _10677_/B _10542_/X _10328_/X _10333_/B vssd1 vssd1 vccd1 vccd1 _10544_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13263_ _13287_/A _13263_/B vssd1 vssd1 vccd1 vccd1 _15107_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10475_ _11542_/A _11606_/A _11536_/A _11168_/A vssd1 vssd1 vccd1 vccd1 _10477_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15002_ _15258_/CLK hold142/X vssd1 vssd1 vccd1 vccd1 _15002_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08033__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12904__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ _12247_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12214_/Y sky130_fd_sc_hd__nor2_1
X_13194_ _13404_/A _13194_/B vssd1 vssd1 vccd1 vccd1 _15059_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output169_A _15181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08584__A2 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ hold2653/X _12173_/A2 _12144_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11918__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12076_ _14978_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12668__A1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10679__B1 _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ _11027_/A _11027_/B _11014_/Y vssd1 vssd1 vccd1 vccd1 _11027_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_0_95_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07416__B _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10123__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10143__A2 _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15263_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_205_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11653__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13093__A1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ hold2765/X _13103_/A2 _13078_/B1 _13198_/B vssd1 vssd1 vccd1 vccd1 _12978_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13153__B _13153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14717_ _15261_/CLK _14717_/D vssd1 vssd1 vccd1 vccd1 _14717_/Q sky130_fd_sc_hd__dfxtp_1
X_11929_ _13651_/A1 hold2253/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11929_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10851__B1 _10850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14648_ _15385_/CLK hold482/X vssd1 vssd1 vccd1 vccd1 hold481/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_28 _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12484__S _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2284_A _13477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _15013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ _15380_/CLK hold206/X vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07120_ _13721_/A1 hold1733/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07120_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07578__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07051_ _13656_/A1 hold1489/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07051_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10017__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11828__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput168 _15180_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[15] sky130_fd_sc_hd__buf_12
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput179 _15190_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[25] sky130_fd_sc_hd__buf_12
XFILLER_0_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07953_ _08677_/A _08892_/A _11566_/A _10507_/A vssd1 vssd1 vccd1 vccd1 _08010_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06904_ _06904_/A vssd1 vssd1 vccd1 vccd1 _13240_/A sky130_fd_sc_hd__inv_2
XANTENNA__11129__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__A _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07884_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _07884_/X sky130_fd_sc_hd__and2_2
XFILLER_0_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09623_ hold2600/X _09344_/B _09346_/B vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_207_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12659__S _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13344__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09554_ _09551_/Y _09552_/X _09411_/Y _09413_/X vssd1 vssd1 vccd1 vccd1 _09555_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09827__A2 _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10687__B _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08505_ _08598_/B _08505_/B vssd1 vssd1 vccd1 vccd1 _08507_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _11288_/A1 _13392_/B _09379_/X vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12831__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07933__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ _08434_/Y _08436_/B vssd1 vssd1 vccd1 vccd1 _08437_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ _08877_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _08367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07318_ _07318_/A _11285_/A vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__and2_1
XANTENNA__07488__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08503_/A sky130_fd_sc_hd__and2_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07249_ _09914_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _07299_/B _07302_/B _10077_/B _07297_/Y vssd1 vssd1 vccd1 vccd1 _10601_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09212__B1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08901__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11738__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10191_/A _10191_/B _10191_/C vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__and3_2
XFILLER_0_121_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08971__C1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__B _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout362 _07337_/Y vssd1 vssd1 vccd1 vccd1 _07390_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07236__B _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13950_ _15415_/CLK _13950_/D vssd1 vssd1 vccd1 vccd1 _13950_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout373 _07812_/X vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__clkbuf_8
Xfanout384 _11895_/X vssd1 vssd1 vccd1 vccd1 _11927_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__11322__B2 _13202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 _07677_/Y vssd1 vssd1 vccd1 vccd1 _07693_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_199_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12901_ _12951_/A _12901_/B vssd1 vssd1 vccd1 vccd1 _12902_/C sky130_fd_sc_hd__or2_1
XFILLER_0_198_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13881_ _15444_/CLK _13881_/D vssd1 vssd1 vccd1 vccd1 _13881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13254__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12832_ _13171_/A _12832_/B vssd1 vssd1 vccd1 vccd1 _14961_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09170__C _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11625__A2 _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12763_ _12917_/B1 _12758_/X _12762_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12770_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _15270_/CLK _14502_/D vssd1 vssd1 vccd1 vccd1 _14502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11714_ hold1771/X _13668_/A1 _11728_/S vssd1 vssd1 vccd1 vccd1 _11714_/X sky130_fd_sc_hd__mux2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12694_ _12700_/S0 _12689_/X _12693_/X _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12695_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14433_ _15305_/CLK _14433_/D vssd1 vssd1 vccd1 vccd1 _14433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11645_ _11645_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11645_/X sky130_fd_sc_hd__and2_1
XFILLER_0_154_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11502__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__B1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 dmemresp_rdata[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14364_ _15263_/CLK _14364_/D vssd1 vssd1 vccd1 vccd1 _14364_/Q sky130_fd_sc_hd__dfxtp_1
X_11576_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__xnor2_1
Xinput26 dmemresp_rdata[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
Xinput37 imemresp_data[13] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 imemresp_data[23] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13315_ input145/X fanout5/X fanout3/X input113/X vssd1 vssd1 vccd1 vccd1 _13315_/X
+ sky130_fd_sc_hd__a22o_1
Xinput59 imemresp_data[4] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
X_10527_ _11561_/A _11378_/D _11542_/B _14947_/Q vssd1 vssd1 vccd1 vccd1 _10528_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10118__A _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14295_ _14909_/CLK hold814/X vssd1 vssd1 vccd1 vccd1 hold813/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08006__A1 _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ input140/X fanout6/X fanout4/X input108/X vssd1 vssd1 vccd1 vccd1 _13246_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08006__B2 _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ _11606_/B _10456_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10460_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12433__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10389_ _10389_/A _10560_/A _10389_/C vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__nor3_1
X_13177_ _13386_/A _13177_/B vssd1 vssd1 vccd1 vccd1 _15042_/D sky130_fd_sc_hd__and2_1
XFILLER_0_97_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ _12128_/A _12128_/B _12128_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12128_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__13148__B _13148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12059_ _12059_/A _12059_/B vssd1 vssd1 vccd1 vccd1 _14842_/D sky130_fd_sc_hd__and2_1
XFILLER_0_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__A2 _14959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13164__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12813__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__B _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09270_ _09271_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _09270_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08493__A1 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08493__B2 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08221_ _10507_/A _08776_/B _11550_/A _08776_/A vssd1 vssd1 vccd1 vccd1 _08222_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08152_ _08152_/A _08152_/B _08152_/C vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__nand3_2
XANTENNA__11412__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__A _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12672__S0 _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12227__B _13749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07101__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _13739_/A1 hold2185/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07103_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08083_ _08082_/B _08082_/C _08082_/A vssd1 vssd1 vccd1 vccd1 _08085_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15304_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ hold397/X _13738_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold398/A sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12424__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09536__B _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12975__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12243__A _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A2 _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2701 _14843_/Q vssd1 vssd1 vccd1 vccd1 hold2701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2712 _14832_/Q vssd1 vssd1 vccd1 vccd1 hold2712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2723 _12056_/X vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08985_ _09941_/A _08985_/B vssd1 vssd1 vccd1 vccd1 _08985_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout484_A _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2734 _13428_/B vssd1 vssd1 vccd1 vccd1 _12271_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2745 _15174_/Q vssd1 vssd1 vccd1 vccd1 hold2745/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _08760_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07936_/Y sky130_fd_sc_hd__nor2_1
Xhold2756 _15169_/Q vssd1 vssd1 vccd1 vccd1 hold2756/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2767 _15110_/Q vssd1 vssd1 vccd1 vccd1 hold2767/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10107__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2778 _09342_/X vssd1 vssd1 vccd1 vccd1 _13391_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07771__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2789 _15103_/Q vssd1 vssd1 vccd1 vccd1 hold2789/X sky130_fd_sc_hd__buf_1
XANTENNA_fanout651_A _15197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ _14100_/Q _14101_/Q _07866_/X _14084_/Q vssd1 vssd1 vccd1 vccd1 _07867_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10698__A _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09606_ _09421_/Y _09461_/A _09604_/Y _09605_/X vssd1 vssd1 vccd1 vccd1 _09606_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07798_ hold475/X _13736_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold476/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09537_ _09537_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12804__A1 _13393_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _09323_/Y _09328_/B _09466_/X _09467_/Y vssd1 vssd1 vccd1 vccd1 _09471_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09108__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08419_ _08512_/B _08418_/B _08418_/C vssd1 vssd1 vccd1 vccd1 _08420_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09399_ _09260_/A _09259_/B _09257_/X vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11430_ _11430_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _11431_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_191_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _11524_/A _11359_/Y _11250_/B _11252_/B vssd1 vssd1 vccd1 vccd1 _11361_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10312_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11791__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ _13096_/X _13097_/X _13099_/X _13098_/X _13100_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _13101_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14080_ _15348_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 _14080_/Q sky130_fd_sc_hd__dfxtp_1
X_11292_ _11290_/Y _11481_/B vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_132_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08539__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13031_ _07355_/Y _13168_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _13032_/B sky130_fd_sc_hd__o21a_1
X_10243_ _14805_/Q _14517_/Q hold919/A _14741_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10244_/B sky130_fd_sc_hd__mux4_1
XANTENNA__07747__A0 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__D _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A1 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _10175_/B vssd1 vssd1 vccd1 vccd1 _10174_/Y sky130_fd_sc_hd__inv_2
X_14982_ _14992_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 _14982_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07681__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13933_ _15042_/CLK _13933_/D vssd1 vssd1 vccd1 vccd1 _13933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13864_ _14783_/CLK _13864_/D vssd1 vssd1 vccd1 vccd1 _13864_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11059__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ hold643/X hold941/X _12915_/S vssd1 vssd1 vccd1 vccd1 _12815_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13795_ _09344_/A _13797_/A2 _13630_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15424_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11931__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08475__A1 _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12746_ hold373/A _15278_/Q hold347/A _14379_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12746_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12677_ _13027_/A _12677_/B _12677_/C vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__and3_1
XFILLER_0_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11232__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14416_ _15062_/CLK hold502/X vssd1 vssd1 vccd1 vccd1 hold501/A sky130_fd_sc_hd__dfxtp_1
X_11628_ _11628_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15396_ _15433_/CLK hold642/X vssd1 vssd1 vccd1 vccd1 hold641/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10034__A1 _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ _15056_/CLK _14347_/D vssd1 vssd1 vccd1 vccd1 _14347_/Q sky130_fd_sc_hd__dfxtp_1
X_11559_ _11566_/A _15225_/Q _11336_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11635_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold607 hold607/A vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 hold618/A vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold629 hold629/A vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14278_ _14731_/CLK hold612/X vssd1 vssd1 vccd1 vccd1 hold611/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13159__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ hold741/X _13675_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold742/A sky130_fd_sc_hd__mux2_1
XANTENNA__12063__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12731__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07833__S0 _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 _11737_/X vssd1 vssd1 vccd1 vccd1 _14531_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2019 _13941_/Q vssd1 vssd1 vccd1 vccd1 hold2019/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 _14798_/Q vssd1 vssd1 vccd1 vccd1 hold1307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08770_ _08755_/Y _08760_/Y _08769_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08771_/B sky130_fd_sc_hd__a221o_1
Xhold1318 _11772_/X vssd1 vssd1 vccd1 vccd1 _14597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07591__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1329 _13812_/Q vssd1 vssd1 vccd1 vccd1 hold1329/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09372__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ hold319/X _13727_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__mux2_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11407__A _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12002__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ hold2039/X _15044_/Q _07660_/S vssd1 vssd1 vccd1 vccd1 _07652_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _13689_/A1 hold1695/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07583_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11841__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ _09321_/B _09321_/C _09321_/A vssd1 vssd1 vccd1 vccd1 _09324_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08138__D _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08466__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09253_ _09253_/A _09435_/A _09714_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09255_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_157_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ _08564_/A1 _08197_/Y _08199_/Y _08201_/Y _08203_/Y vssd1 vssd1 vccd1 vccd1
+ _08204_/X sky130_fd_sc_hd__o32a_1
X_09184_ _09184_/A _09184_/B _09184_/C vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ hold2516/X input29/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13178_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07766__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _15395_/Q _14530_/Q _14690_/Q _14754_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08066_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_114_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07017_ hold809/X _13655_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 hold810/A sky130_fd_sc_hd__mux2_1
XANTENNA__12948__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2520 _07389_/Y vssd1 vssd1 vccd1 vccd1 hold2520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2531 _15144_/Q vssd1 vssd1 vccd1 vccd1 hold2531/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2542 _15002_/Q vssd1 vssd1 vccd1 vccd1 hold2542/X sky130_fd_sc_hd__buf_2
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _08852_/B _08854_/B _08850_/X vssd1 vssd1 vccd1 vccd1 _08969_/B sky130_fd_sc_hd__a21o_1
Xhold2553 _14995_/Q vssd1 vssd1 vccd1 vccd1 hold2553/X sky130_fd_sc_hd__buf_2
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2564 _15001_/Q vssd1 vssd1 vccd1 vccd1 hold2564/X sky130_fd_sc_hd__buf_2
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2575 _15338_/Q vssd1 vssd1 vccd1 vccd1 _07346_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1830 _07758_/X vssd1 vssd1 vccd1 vccd1 _14374_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2586 _14976_/Q vssd1 vssd1 vccd1 vccd1 hold2586/X sky130_fd_sc_hd__buf_2
Xhold1841 _14499_/Q vssd1 vssd1 vccd1 vccd1 hold1841/X sky130_fd_sc_hd__dlygate4sd3_1
X_07919_ _07919_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07920_/B sky130_fd_sc_hd__nand2_1
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1852 _07489_/X vssd1 vssd1 vccd1 vccd1 _14117_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2597 _11300_/X vssd1 vssd1 vccd1 vccd1 _14453_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08899_ _08897_/X _08899_/B vssd1 vssd1 vccd1 vccd1 _08900_/B sky130_fd_sc_hd__and2b_1
Xhold1863 _14127_/Q vssd1 vssd1 vccd1 vccd1 hold1863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1874 _07175_/X vssd1 vssd1 vccd1 vccd1 _13983_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1885 _15267_/Q vssd1 vssd1 vccd1 vccd1 hold1885/X sky130_fd_sc_hd__dlygate4sd3_1
X_10930_ _13890_/Q hold293/A _13858_/Q _13826_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10930_/X sky130_fd_sc_hd__mux4_1
Xhold1896 _11761_/X vssd1 vssd1 vccd1 vccd1 _14555_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07006__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10861_ _11550_/A _11620_/B _15221_/Q _11526_/A vssd1 vssd1 vccd1 vccd1 _10863_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11751__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12596_/X _12597_/X _12599_/X _12598_/X _12644_/A1 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12601_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_112_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13580_ _13580_/A _13586_/B vssd1 vssd1 vccd1 vccd1 _13580_/Y sky130_fd_sc_hd__nand2_1
X_10792_ _10792_/A _10792_/B vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09654__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _08345_/A _08636_/A _13148_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12532_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08552__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15250_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12462_ _12689_/S1 _12459_/X _12461_/X vssd1 vssd1 vccd1 vccd1 _12462_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10016__A1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201_ _15087_/CLK _14201_/D vssd1 vssd1 vccd1 vccd1 _14201_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13678__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__A1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10016__B2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11413_ _11569_/A _11605_/B _11414_/C _11608_/A vssd1 vssd1 vccd1 vccd1 _11416_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09501__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _15188_/CLK _15181_/D vssd1 vssd1 vccd1 vccd1 _15181_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12393_ _12599_/S1 _12390_/X _12392_/X vssd1 vssd1 vccd1 vccd1 _12393_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10567__A2 _10566_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__C _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12961__B1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ _14775_/CLK _14132_/D vssd1 vssd1 vccd1 vccd1 _14132_/Q sky130_fd_sc_hd__dfxtp_1
X_11344_ _11344_/A _11344_/B vssd1 vssd1 vccd1 vccd1 _11346_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08361__A _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14063_ _15425_/CLK _14063_/D vssd1 vssd1 vccd1 vccd1 _14063_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12939__S1 _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ _11468_/A _11273_/Y _11051_/X _11054_/Y vssd1 vssd1 vccd1 vccd1 _11276_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13014_ hold599/X hold835/X hold493/X hold999/X _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13014_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10226_ _10221_/X _10222_/X _10225_/Y vssd1 vssd1 vccd1 vccd1 _13397_/B sky130_fd_sc_hd__a21o_4
XANTENNA_output249_A _14453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _10156_/B _10156_/C _10156_/A vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_14965_ _14971_/CLK _14965_/D vssd1 vssd1 vccd1 vccd1 _14965_/Q sky130_fd_sc_hd__dfxtp_1
X_10088_ _10426_/A _10087_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _10088_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_169_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13916_ _15449_/CLK _13916_/D vssd1 vssd1 vccd1 vccd1 _13916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10131__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14896_ _14989_/CLK _14896_/D vssd1 vssd1 vccd1 vccd1 _14896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ _15276_/CLK _13847_/D vssd1 vssd1 vccd1 vccd1 _13847_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11661__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13778_ hold205/X vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12875__S0 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10255__A1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13161__B _13161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12729_ _09209_/Y _13104_/A2 _12728_/X vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15448_ _15448_/CLK _15448_/D vssd1 vssd1 vccd1 vccd1 _15448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15379_ _15379_/CLK hold448/X vssd1 vssd1 vccd1 vccd1 hold447/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07586__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 hold404/A vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold415 hold415/A vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold426 hold426/A vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 hold437/A vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08702__C _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold448 hold448/A vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold459 hold459/A vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09940_ hold793/A _14515_/Q _14643_/Q _14739_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09941_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09871_ _09871_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09872_/B sky130_fd_sc_hd__nor2_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11836__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _08710_/Y _08714_/B _08820_/Y _08821_/X vssd1 vssd1 vccd1 vccd1 _08825_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__08923__A2 _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1104 _11965_/X vssd1 vssd1 vccd1 vccd1 _14784_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 _14154_/Q vssd1 vssd1 vccd1 vccd1 hold1115/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _07694_/X vssd1 vssd1 vccd1 vccd1 _14314_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _14757_/Q vssd1 vssd1 vccd1 vccd1 hold1137/X sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ _13875_/Q _14003_/Q _13843_/Q _13811_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08753_/X sky130_fd_sc_hd__mux4_1
Xhold1148 _07214_/X vssd1 vssd1 vccd1 vccd1 _14021_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _14765_/Q vssd1 vssd1 vccd1 vccd1 hold1159/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ hold961/X hold2765/A _07709_/S vssd1 vssd1 vccd1 vccd1 hold962/A sky130_fd_sc_hd__mux2_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _09026_/B _08685_/C _09712_/A _08908_/A vssd1 vssd1 vccd1 vccd1 _08686_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13680__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07635_ hold1295/X _13741_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07635_/X sky130_fd_sc_hd__mux2_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout447_A _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13352__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ _13396_/A hold209/X vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__and2_1
XANTENNA__08439__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__A1 _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _09305_/A _09305_/B _09305_/C vssd1 vssd1 vccd1 vccd1 _09307_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07350__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout614_A _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07497_ hold1747/X _13736_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07497_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09236_ _09514_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09236_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09167_ _09167_/A _09167_/B vssd1 vssd1 vccd1 vccd1 _09175_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_161_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__S _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07496__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09277__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _08869_/A _08115_/X _08117_/X vssd1 vssd1 vccd1 vccd1 _08118_/Y sky130_fd_sc_hd__o21ai_1
X_09098_ _09941_/A _09095_/X _09097_/X vssd1 vssd1 vccd1 vccd1 _09098_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09708__C _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _13546_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08049_/Y sky130_fd_sc_hd__nor2_1
Xhold960 hold960/A vssd1 vssd1 vccd1 vccd1 hold960/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold971 hold971/A vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _11541_/A _11351_/B _11614_/B _11586_/B vssd1 vssd1 vccd1 vccd1 _11242_/A
+ sky130_fd_sc_hd__nand4_2
Xhold982 hold982/A vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 hold993/A vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _10011_/A _10011_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__or2_1
XANTENNA__11746__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__A1 hold2593/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2350 _14061_/Q vssd1 vssd1 vccd1 vccd1 _06920_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2361 _12179_/X vssd1 vssd1 vccd1 vccd1 _14900_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2372 _15041_/Q vssd1 vssd1 vccd1 vccd1 hold2372/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2383 _13551_/X vssd1 vssd1 vccd1 vccd1 _15301_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2394 _15004_/Q vssd1 vssd1 vccd1 vccd1 _12128_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1660 _13711_/X vssd1 vssd1 vccd1 vccd1 _15417_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07244__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14750_/CLK _14750_/D vssd1 vssd1 vccd1 vccd1 _14750_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1671 _14128_/Q vssd1 vssd1 vccd1 vccd1 hold1671/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1682 _07096_/X vssd1 vssd1 vccd1 vccd1 _13909_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11962_ hold589/X _13651_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 hold590/A sky130_fd_sc_hd__mux2_1
XANTENNA__09875__B1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1693 _14123_/Q vssd1 vssd1 vccd1 vccd1 hold1693/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__A0 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ hold1221/X _13734_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 _13701_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _10958_/A _10737_/X _10734_/A vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__o21ai_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _15455_/CLK hold652/X vssd1 vssd1 vccd1 vccd1 hold651/A sky130_fd_sc_hd__dfxtp_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ hold655/X _13714_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold656/A sky130_fd_sc_hd__mux2_1
XFILLER_0_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ input42/X _13634_/B vssd1 vssd1 vccd1 vccd1 _13632_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10844_ _10844_/A _10844_/B _10844_/C vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12226__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07260__A _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13563_ _08851_/A _09222_/B _13562_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _13563_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ _10760_/Y _10765_/Y _10774_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _10776_/B sky130_fd_sc_hd__a221o_1
XANTENNA__08075__B _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15302_ _15304_/CLK _15302_/D vssd1 vssd1 vccd1 vccd1 _15302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ hold379/A hold495/A _14146_/Q _14464_/Q _12566_/S _12368_/A vssd1 vssd1 vccd1
+ vccd1 _12514_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_125_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08850__A1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ _13499_/A hold41/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__and2_1
XFILLER_0_164_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15233_ _15250_/CLK _15233_/D vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12445_ _12445_/A _12445_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08803__B _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__A1 _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ _15325_/CLK _15164_/D vssd1 vssd1 vccd1 vccd1 _15164_/Q sky130_fd_sc_hd__dfxtp_1
X_12376_ _12669_/A1 _12371_/X _12375_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12376_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08602__B2 _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12325__B _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ _15436_/CLK _14115_/D vssd1 vssd1 vccd1 vccd1 _14115_/Q sky130_fd_sc_hd__dfxtp_1
X_11327_ _11236_/A _11236_/B _11238_/X vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10126__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07419__B _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ _15384_/CLK hold524/X vssd1 vssd1 vccd1 vccd1 hold523/A sky130_fd_sc_hd__dfxtp_1
X_14046_ _14105_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dfxtp_1
X_11258_ _11258_/A _11329_/A _11258_/C vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11656__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10209_ _10206_/X _10207_/Y _10053_/Y _10055_/X vssd1 vssd1 vccd1 vccd1 _10209_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13437__A _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12341__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11189_ _11586_/A _11614_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _11189_/X sky130_fd_sc_hd__and3_1
XANTENNA__08461__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13156__B _13156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _15225_/CLK _14948_/D vssd1 vssd1 vccd1 vccd1 _14948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08669__B2 _13184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ _14987_/CLK _14879_/D vssd1 vssd1 vccd1 vccd1 _14879_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13172__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07420_ hold195/X _07475_/B vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__and2_1
XFILLER_0_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12848__S0 _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07351_ _07351_/A _07351_/B _07360_/B _07351_/D vssd1 vssd1 vccd1 vccd1 _07359_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_58_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A2 _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07282_ _08012_/B _10507_/A vssd1 vssd1 vccd1 vccd1 _07283_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09021_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _09021_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2746_A _15175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11728__A1 _15068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10087__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10936__C1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10400__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13025__S0 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _14445_/Q _09923_/B vssd1 vssd1 vccd1 vccd1 _10082_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 hold285/X vssd1 vssd1 vccd1 vccd1 _13659_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout714 _13719_/A1 vssd1 vssd1 vccd1 vccd1 _13653_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12153__A1 hold2617/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 _14961_/Q vssd1 vssd1 vccd1 vccd1 _11605_/B sky130_fd_sc_hd__buf_6
XANTENNA_fanout397_A _07610_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 _11390_/A vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13347__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09856_/B sky130_fd_sc_hd__xnor2_2
Xfanout747 _14952_/Q vssd1 vssd1 vccd1 vccd1 _11564_/A sky130_fd_sc_hd__buf_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout758 _11620_/A vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__buf_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout769 _08926_/A vssd1 vssd1 vccd1 vccd1 _10185_/A sky130_fd_sc_hd__buf_6
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__nand2_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09780_/A _13586_/B _09784_/Y _13579_/C1 vssd1 vssd1 vccd1 vccd1 _09785_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout564_A _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ _13669_/A1 hold1801/X _07010_/S vssd1 vssd1 vccd1 vccd1 _06997_/X sky130_fd_sc_hd__mux2_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _10024_/A _08570_/Y _07320_/B vssd1 vssd1 vccd1 vccd1 _08846_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09857__B1 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_107 hold2653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout731_A _14958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_129 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _12252_/B _08667_/B vssd1 vssd1 vccd1 vccd1 _08667_/Y sky130_fd_sc_hd__nor2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout829_A _14488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07618_ hold1367/X _13724_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07618_/X sky130_fd_sc_hd__mux2_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08598_/A _08598_/B vssd1 vssd1 vccd1 vccd1 _08612_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12839__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07549_ _13386_/A hold233/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__and2_1
XANTENNA__12613__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_87_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07096__A0 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _10560_/A _10560_/B _10560_/C vssd1 vssd1 vccd1 vccd1 _10561_/B sky130_fd_sc_hd__or3_1
XFILLER_0_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clk_A clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09219_ _15149_/Q _09925_/A2 _09494_/A1 vssd1 vssd1 vccd1 vccd1 _09219_/Y sky130_fd_sc_hd__a21oi_1
X_10491_ _10491_/A _10491_/B _10491_/C vssd1 vssd1 vccd1 vccd1 _10494_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12426__A _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ hold755/A _13799_/Q _12237_/S vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11195__A2 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12392__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09793__C1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__B _14970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ hold2562/X _12173_/A2 _12160_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12161_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12860__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_145_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ _11112_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _13370_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12092_ _14986_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12092_/X
+ sky130_fd_sc_hd__or4_1
Xhold790 hold790/A vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08348__B1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13257__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ _11566_/A _15223_/Q _11229_/A _11042_/D vssd1 vssd1 vccd1 vccd1 _11045_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10155__B1 _10154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13691__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2180 _07058_/X vssd1 vssd1 vccd1 vccd1 _13874_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2191 _14036_/Q vssd1 vssd1 vccd1 vccd1 _07461_/A sky130_fd_sc_hd__dlygate4sd3_1
X_14802_ _15379_/CLK _14802_/D vssd1 vssd1 vccd1 vccd1 _14802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _13050_/S0 _12989_/X _12993_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _12995_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10458__A1 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1490 _07051_/X vssd1 vssd1 vccd1 vccd1 _13867_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _15190_/CLK _14733_/D vssd1 vssd1 vccd1 vccd1 _14733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11945_ _13700_/A1 hold1159/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11945_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _15438_/CLK _14664_/D vssd1 vssd1 vccd1 vccd1 _14664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ hold1755/X _13730_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11876_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13615_ input64/X _13636_/B vssd1 vssd1 vccd1 vccd1 _13615_/X sky130_fd_sc_hd__or2_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10827_ _14953_/Q _11536_/A _10827_/C _10827_/D vssd1 vssd1 vccd1 vccd1 _10830_/C
+ sky130_fd_sc_hd__nand4_1
X_14595_ _14595_/CLK _14595_/D vssd1 vssd1 vccd1 vccd1 _14595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13546_ _13546_/A _13554_/B vssd1 vssd1 vccd1 vccd1 _13546_/X sky130_fd_sc_hd__or2_1
XANTENNA__08284__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ _13889_/Q hold775/A _13857_/Q _13825_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10758_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_171_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _13477_/A _13477_/B vssd1 vssd1 vccd1 vccd1 _13477_/X sky130_fd_sc_hd__and2_1
X_10689_ _10515_/B _10517_/B _10515_/A vssd1 vssd1 vccd1 vccd1 _10691_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_113_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15216_ _15222_/CLK _15216_/D vssd1 vssd1 vccd1 vccd1 _15216_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09379__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ hold2372/X _12329_/B _12953_/B1 _13176_/B vssd1 vssd1 vccd1 vccd1 _12428_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput306 _14867_/Q vssd1 vssd1 vccd1 vccd1 out1[22] sky130_fd_sc_hd__buf_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput317 _14848_/Q vssd1 vssd1 vccd1 vccd1 out1[3] sky130_fd_sc_hd__buf_12
Xoutput328 _14826_/Q vssd1 vssd1 vccd1 vccd1 out2[13] sky130_fd_sc_hd__buf_12
XFILLER_0_140_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15147_ _15309_/CLK _15147_/D vssd1 vssd1 vccd1 vccd1 _15147_/Q sky130_fd_sc_hd__dfxtp_1
X_12359_ _12607_/A _12359_/B vssd1 vssd1 vccd1 vccd1 _14942_/D sky130_fd_sc_hd__nor2_1
Xoutput339 _14836_/Q vssd1 vssd1 vccd1 vccd1 out2[23] sky130_fd_sc_hd__buf_12
XFILLER_0_168_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09645__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _15270_/CLK hold890/X vssd1 vssd1 vccd1 vccd1 hold889/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12135__A1 _12068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ _14083_/CLK _14029_/D vssd1 vssd1 vccd1 vccd1 _14029_/Q sky130_fd_sc_hd__dfxtp_1
X_06920_ _06920_/A vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__inv_2
XANTENNA__13167__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10697__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__B2 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__B _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09570_ _09571_/A _09714_/A _09714_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09570_/X
+ sky130_fd_sc_hd__and4_1
X_08521_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08521_/X sky130_fd_sc_hd__xor2_1
XANTENNA__10449__A1 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2696_A _14844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__B2 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09811__C _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08452_ _12243_/A _08452_/B vssd1 vssd1 vccd1 vccd1 _08452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07403_ _07403_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14033_/D sky130_fd_sc_hd__nor2_1
X_08383_ _09860_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13630__A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07334_ hold2820/X _08849_/A _07334_/C _07334_/D vssd1 vssd1 vccd1 vccd1 _07359_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ _11605_/A _10306_/A vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_27_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09004_ _09435_/A _09571_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _09004_/X sky130_fd_sc_hd__and3_1
XFILLER_0_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ hold1971/X _13664_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07196_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12374__A1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07774__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout500 _06943_/Y vssd1 vssd1 vccd1 vccd1 _13100_/S0 sky130_fd_sc_hd__buf_8
XANTENNA_fanout779_A _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _10252_/A vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__buf_6
X_09906_ _09903_/A _09904_/X _09667_/Y _09670_/Y vssd1 vssd1 vccd1 vccd1 _09906_/Y
+ sky130_fd_sc_hd__o211ai_2
Xfanout522 _08880_/A1 vssd1 vssd1 vccd1 vccd1 _08992_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__13077__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout533 _15424_/Q vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__clkbuf_8
Xfanout544 _12211_/S1 vssd1 vssd1 vccd1 vccd1 _12244_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout555 _11501_/S1 vssd1 vssd1 vccd1 vccd1 _11506_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout566 _10087_/S0 vssd1 vssd1 vccd1 vccd1 _09239_/S0 sky130_fd_sc_hd__buf_8
X_09837_ _09684_/Y _09686_/X _09835_/Y _09836_/X vssd1 vssd1 vccd1 vccd1 _09839_/B
+ sky130_fd_sc_hd__a211oi_2
Xfanout577 _07448_/A vssd1 vssd1 vccd1 vccd1 _10744_/A sky130_fd_sc_hd__buf_4
Xfanout588 _15215_/Q vssd1 vssd1 vccd1 vccd1 _11536_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__08976__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 _09676_/D vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__buf_4
X_09768_ _09767_/B _09767_/C _09767_/A vssd1 vssd1 vccd1 vccd1 _09914_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12429__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08719_ _08611_/Y _08613_/X _08716_/X _08718_/Y vssd1 vssd1 vccd1 vccd1 _08721_/B
+ sky130_fd_sc_hd__a211o_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _10002_/C _10283_/C _10115_/D _09846_/B vssd1 vssd1 vccd1 vccd1 _09702_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11730_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _11762_/S sky130_fd_sc_hd__or2_4
XFILLER_0_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07014__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ _13725_/A1 hold1567/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ _13481_/A _13400_/B vssd1 vssd1 vccd1 vccd1 _15191_/D sky130_fd_sc_hd__and2_1
XFILLER_0_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12062__A0 _12128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ _10612_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10614_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14380_ _15376_/CLK _14380_/D vssd1 vssd1 vccd1 vccd1 _14380_/Q sky130_fd_sc_hd__dfxtp_1
X_11592_ _11592_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _11602_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ input86/X fanout2/X _13330_/X vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10543_ _10328_/X _10333_/B _10677_/B _10542_/X vssd1 vssd1 vccd1 vccd1 _10543_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11060__A _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13262_ input93/X fanout1/X _13261_/X vssd1 vssd1 vccd1 vccd1 _13263_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _11168_/A _11542_/A _11606_/A _11536_/A vssd1 vssd1 vccd1 vccd1 _10477_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15001_ _15258_/CLK hold102/X vssd1 vssd1 vccd1 vccd1 _15001_/Q sky130_fd_sc_hd__dfxtp_1
X_12213_ _14653_/Q _13926_/Q _15427_/Q _13894_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12214_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13686__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12590__S _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ _13397_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _15058_/D sky130_fd_sc_hd__and2_1
XANTENNA__08033__A2 _13378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07684__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _14883_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09518__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12075_ hold2452/X _12099_/A2 _12074_/X _13492_/A vssd1 vssd1 vccd1 vccd1 _12075_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10404__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10679__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _11025_/A _11025_/B _11025_/C vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10679__B2 _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10123__B _14964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11934__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2__f_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__B _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13434__B _13434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _13102_/A _12977_/B _12977_/C vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__and3_1
XFILLER_0_204_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ _15455_/CLK hold572/X vssd1 vssd1 vccd1 vccd1 hold571/A sky130_fd_sc_hd__dfxtp_1
X_11928_ _11928_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _11960_/S sky130_fd_sc_hd__or2_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14647_ _15191_/CLK _14647_/D vssd1 vssd1 vccd1 vccd1 _14647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12765__S _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ hold877/X _13746_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold878/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14578_ _15379_/CLK hold202/X vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_29 _14923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13529_ hold2765/A hold449/X _13534_/S vssd1 vssd1 vccd1 vccd1 hold450/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12066__A _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07050_ _13655_/A1 hold1751/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07050_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_180_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12356__A1 _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10017__C _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput169 _15181_/Q vssd1 vssd1 vccd1 vccd1 dmemreq_addr[16] sky130_fd_sc_hd__buf_12
XFILLER_0_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07952_ _08892_/A _11566_/A _10507_/A _08677_/A vssd1 vssd1 vccd1 vccd1 _07952_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__10314__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06903_ _06903_/A vssd1 vssd1 vccd1 vccd1 _12294_/A sky130_fd_sc_hd__inv_2
X_07883_ hold2694/X input23/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13174_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_207_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10033__B _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ _11288_/A1 _13393_/B _09521_/X vssd1 vssd1 vccd1 vccd1 _13444_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13069__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ _09411_/Y _09413_/X _09551_/Y _09552_/X vssd1 vssd1 vccd1 vccd1 _09555_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_195_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08504_ _08598_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08505_/B sky130_fd_sc_hd__nand2_1
X_09484_ _09615_/B _09479_/X _09483_/X vssd1 vssd1 vccd1 vccd1 _13392_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12831__A2 _13160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout527_A _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__A0 hold2553/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13360__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07769__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ _14275_/Q hold577/A _14147_/Q _14465_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08367_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08454__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07317_ _15225_/Q _14969_/Q vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _11564_/B _11605_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__or2_1
XFILLER_0_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07179_ _13746_/A1 hold1931/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07179_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08901__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _10189_/B _10189_/C _10189_/A vssd1 vssd1 vccd1 vccd1 _10191_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13238__C _15355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07009__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout363 _13027_/A vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__buf_6
Xfanout374 _07812_/X vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11322__A2 _07899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 _11745_/S vssd1 vssd1 vccd1 vccd1 _11761_/S sky130_fd_sc_hd__clkbuf_16
X_12900_ _12896_/X _12897_/X _12899_/X _12898_/X _12950_/S0 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12901_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11754__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _07677_/Y vssd1 vssd1 vccd1 vccd1 _07709_/S sky130_fd_sc_hd__clkbuf_16
X_13880_ _15087_/CLK _13880_/D vssd1 vssd1 vccd1 vccd1 _13880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _13106_/A1 _13160_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12832_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12949_/S1 _12759_/X _12761_/X vssd1 vssd1 vccd1 vccd1 _12762_/X sky130_fd_sc_hd__a21o_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__D _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _15400_/CLK hold710/X vssd1 vssd1 vccd1 vccd1 hold709/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ hold1413/X _13519_/A0 _11728_/S vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__mux2_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12585__S _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12693_ _12699_/S1 _12690_/X _12692_/X vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__a21o_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07679__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14432_ _15305_/CLK _14432_/D vssd1 vssd1 vccd1 vccd1 _14432_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_166_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11644_ _11645_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11644_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12586__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ _15364_/CLK _14363_/D vssd1 vssd1 vccd1 vccd1 _14363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11575_ _11575_/A _11575_/B vssd1 vssd1 vccd1 vccd1 _11576_/B sky130_fd_sc_hd__xnor2_1
Xinput16 dmemresp_rdata[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput27 dmemresp_rdata[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
XFILLER_0_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13314_ _13317_/A _13314_/B vssd1 vssd1 vccd1 vccd1 _15124_/D sky130_fd_sc_hd__nor2_1
Xinput38 imemresp_data[14] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_1
XFILLER_0_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput49 imemresp_data[24] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10526_ _11541_/A _11351_/B _11378_/D _11542_/B vssd1 vssd1 vccd1 vccd1 _10696_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_134_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ _14485_/CLK hold600/X vssd1 vssd1 vccd1 vccd1 hold599/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output181_A _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11929__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ _13287_/A _13245_/B vssd1 vssd1 vccd1 vccd1 _15101_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_150_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08006__A2 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10457_ _11573_/A _11606_/B _11570_/B _11590_/A vssd1 vssd1 vccd1 vccd1 _10457_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12433__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ _13477_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _15041_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10388_ _10387_/A _10387_/B _10387_/C vssd1 vssd1 vccd1 vccd1 _10389_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12127_ hold2483/X _12129_/A2 _12126_/X _12063_/A vssd1 vssd1 vccd1 vccd1 _12127_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07427__B _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ hold2542/X hold2713/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12059_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_165_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11664__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _11564_/A _11378_/C _11010_/C _11010_/D vssd1 vssd1 vccd1 vccd1 _11009_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_205_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08190__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__A _08179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13164__B _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08493__A2 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _08776_/A _10507_/A _08776_/B _11550_/A vssd1 vssd1 vccd1 vccd1 _08222_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12026__A0 hold2538/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13180__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08274__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ _08082_/A _08082_/C _08082_/B vssd1 vssd1 vccd1 vccd1 _08152_/C sky130_fd_sc_hd__o21bai_2
XFILLER_0_133_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11412__B _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08876__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12672__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07102_ _13738_/A1 hold1699/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07102_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08082_ _08082_/A _08082_/B _08082_/C vssd1 vssd1 vccd1 vccd1 _08085_/A sky130_fd_sc_hd__or3_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11839__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07033_ hold659/X _13671_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold660/A sky130_fd_sc_hd__mux2_1
XFILLER_0_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12424__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10044__A _10044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2702 _12060_/X vssd1 vssd1 vccd1 vccd1 _12061_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08984_ hold463/A hold601/A hold747/A hold857/A _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _08985_/B sky130_fd_sc_hd__mux4_1
Xhold2713 _14842_/Q vssd1 vssd1 vccd1 vccd1 hold2713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2724 _14826_/Q vssd1 vssd1 vccd1 vccd1 hold2724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2735 _15057_/Q vssd1 vssd1 vccd1 vccd1 hold2735/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ _08201_/A _07932_/X _07934_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _07936_/B
+ sky130_fd_sc_hd__o211a_1
Xhold2746 _15175_/Q vssd1 vssd1 vccd1 vccd1 hold2746/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2757 _15101_/Q vssd1 vssd1 vccd1 vccd1 hold2757/X sky130_fd_sc_hd__buf_1
XANTENNA_fanout477_A _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2768 _15194_/Q vssd1 vssd1 vccd1 vccd1 hold2768/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2779 _15130_/Q vssd1 vssd1 vccd1 vccd1 hold2779/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__13355__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07866_ _14102_/Q _14104_/Q _14103_/Q _14105_/Q vssd1 vssd1 vccd1 vccd1 _07866_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10698__B _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09605_ _09601_/X _09603_/Y _09461_/C _09464_/B vssd1 vssd1 vccd1 vccd1 _09605_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout644_A _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ hold583/X _13735_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold584/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09536_ _10351_/A _10166_/C vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_211_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08883__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12804__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09130__B1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12360__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09463_/X _09465_/Y _09317_/X _09321_/B vssd1 vssd1 vccd1 vccd1 _09467_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_210_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout811_A _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07499__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08418_ _08512_/B _08418_/B _08418_/C vssd1 vssd1 vccd1 vccd1 _08516_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11603__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _09398_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12568__A1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08349_ _09918_/A _12268_/B _13350_/B _08256_/A _08348_/Y vssd1 vssd1 vccd1 vccd1
+ _08349_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09433__A1 _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08867__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11250_/B _11252_/B _11524_/A _11359_/Y vssd1 vssd1 vccd1 vccd1 _11524_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10311_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11749__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11291_ _11645_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11481_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08631__B _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13080_/A1 _13029_/X hold2776/X vssd1 vssd1 vccd1 vccd1 _13168_/B sky130_fd_sc_hd__a21oi_2
X_10242_ hold843/A hold625/A hold741/A _14386_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10242_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11543__A2 _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _14942_/Q _11586_/B vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07247__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14981_ _15251_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _14981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ _14754_/CLK _13932_/D vssd1 vssd1 vccd1 vccd1 _13932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__A _15227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13863_ _15427_/CLK _13863_/D vssd1 vssd1 vccd1 vccd1 _13863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11059__A1 _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ hold805/X _14222_/Q hold515/X hold1763/X _12841_/S _06942_/A vssd1 vssd1
+ vccd1 vccd1 _12814_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_202_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__B2 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ hold2331/X _13797_/A2 _13628_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _13794_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10806__A1 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12745_ _12745_/A _12745_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12752_/B sky130_fd_sc_hd__or3b_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08475__A2 _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12008__A0 hold2628/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12676_/A _12676_/B vssd1 vssd1 vccd1 vccd1 _12677_/C sky130_fd_sc_hd__or2_1
XFILLER_0_182_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14415_ _15448_/CLK _14415_/D vssd1 vssd1 vccd1 vccd1 _14415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11232__B _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ _11626_/A _11626_/B _11626_/C vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15395_ _15395_/CLK _15395_/D vssd1 vssd1 vccd1 vccd1 _15395_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10129__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09918__A _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ _15374_/CLK hold540/X vssd1 vssd1 vccd1 vccd1 hold539/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08632__C1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _11558_/A _11558_/B vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11659__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 hold608/A vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10509_ _11566_/A _11620_/B vssd1 vssd1 vccd1 vccd1 _10510_/C sky130_fd_sc_hd__and2_1
XFILLER_0_204_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14277_ _15080_/CLK hold994/X vssd1 vssd1 vccd1 vccd1 hold993/A sky130_fd_sc_hd__dfxtp_1
Xhold619 hold619/A vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ _14454_/Q _11650_/B _11476_/Y hold2329/X _13459_/A vssd1 vssd1 vccd1 vccd1
+ _11489_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_100_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13228_ hold1757/X _13674_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13159__B _13159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12731__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13389_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _15024_/D sky130_fd_sc_hd__nor2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2009 _14745_/Q vssd1 vssd1 vccd1 vccd1 hold2009/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07833__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 _11979_/X vssd1 vssd1 vccd1 vccd1 _14798_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10799__A _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1319 _13973_/Q vssd1 vssd1 vccd1 vccd1 hold1319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13175__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ hold499/X _13693_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold500/A sky130_fd_sc_hd__mux2_1
XANTENNA__09360__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__B _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ hold1559/X _13690_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 _07651_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07582_ _13721_/A1 hold1485/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07582_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09321_ _09321_/A _09321_/B _09321_/C vssd1 vssd1 vccd1 vccd1 _09464_/A sky130_fd_sc_hd__and3_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09252_ _09253_/A _09435_/A _09864_/C _09714_/D vssd1 vssd1 vccd1 vccd1 _09252_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07112__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ _08197_/A _08202_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _08203_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ _09180_/X _09181_/Y _09049_/X _09051_/Y vssd1 vssd1 vccd1 vccd1 _09184_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08134_ _12252_/B _08134_/B vssd1 vssd1 vccd1 vccd1 _08134_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09828__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08065_ _08065_/A _08065_/B vssd1 vssd1 vccd1 vccd1 _08065_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_141_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07348__A _15355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07016_ hold1425/X _13687_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07016_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07729__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_A _15213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07782__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2510 _12163_/X vssd1 vssd1 vccd1 vccd1 _14892_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2521 _15109_/Q vssd1 vssd1 vccd1 vccd1 hold2521/X sky130_fd_sc_hd__buf_1
Xhold2532 _08644_/X vssd1 vssd1 vccd1 vccd1 hold2532/X sky130_fd_sc_hd__dlygate4sd3_1
X_08967_ _08965_/X _08967_/B vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__and2b_1
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2543 _12191_/X vssd1 vssd1 vccd1 vccd1 _14906_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2554 _12177_/X vssd1 vssd1 vccd1 vccd1 _14899_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout859_A _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1820 _07623_/X vssd1 vssd1 vccd1 vccd1 _14246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2565 _12189_/X vssd1 vssd1 vccd1 vccd1 _14905_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__B _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1831 _14237_/Q vssd1 vssd1 vccd1 vccd1 hold1831/X sky130_fd_sc_hd__dlygate4sd3_1
X_07918_ _07919_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07920_/A sky130_fd_sc_hd__or2_1
XANTENNA__12486__B1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2576 _14452_/Q vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ _08895_/Y _08896_/X _08780_/X _08782_/X vssd1 vssd1 vccd1 vccd1 _08899_/B
+ sky130_fd_sc_hd__a211o_1
Xhold2587 _12139_/X vssd1 vssd1 vccd1 vccd1 _14880_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1842 _11703_/X vssd1 vssd1 vccd1 vccd1 _14499_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08179__A _08179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__A1 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1853 _14004_/Q vssd1 vssd1 vccd1 vccd1 hold1853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2598 _14427_/Q vssd1 vssd1 vccd1 vccd1 _08042_/B sky130_fd_sc_hd__buf_1
Xhold1864 _07499_/X vssd1 vssd1 vccd1 vccd1 _14127_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1875 _13914_/Q vssd1 vssd1 vccd1 vccd1 hold1875/X sky130_fd_sc_hd__dlygate4sd3_1
X_07849_ _07848_/X _07849_/B _07856_/B _14056_/Q vssd1 vssd1 vccd1 vccd1 _07849_/X
+ sky130_fd_sc_hd__and4b_1
Xhold1886 _13509_/X vssd1 vssd1 vccd1 vccd1 _15267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1897 _14742_/Q vssd1 vssd1 vccd1 vccd1 hold1897/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07901__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07901__B2 _13174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10860_ _11526_/A _11550_/A _11620_/B _15221_/Q vssd1 vssd1 vccd1 vccd1 _10863_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12238__B1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07811__A _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ _11320_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10791_ _10792_/A _10792_/B vssd1 vssd1 vccd1 vccd1 _10791_/Y sky130_fd_sc_hd__nor2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11333__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ _12327_/A _12529_/X _12527_/X vssd1 vssd1 vccd1 vccd1 _13148_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07022__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ _12642_/A1 _12460_/X _12644_/A1 vssd1 vssd1 vccd1 vccd1 _12461_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _15087_/CLK _14200_/D vssd1 vssd1 vccd1 vccd1 _14200_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10016__A2 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _11594_/A _11563_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _11608_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__09957__A2 _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15180_ _15184_/CLK _15180_/D vssd1 vssd1 vccd1 vccd1 _15180_/Q sky130_fd_sc_hd__dfxtp_2
X_12392_ _12642_/A1 _12391_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12392_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09501__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12961__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__C1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ _14419_/CLK _14131_/D vssd1 vssd1 vccd1 vccd1 _14131_/Q sky130_fd_sc_hd__dfxtp_1
X_11343_ _11343_/A _11343_/B _11343_/C vssd1 vssd1 vccd1 vccd1 _11344_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14062_ _15425_/CLK _14062_/D vssd1 vssd1 vccd1 vccd1 _14062_/Q sky130_fd_sc_hd__dfxtp_1
X_11274_ _11051_/X _11054_/Y _11468_/A _11273_/Y vssd1 vssd1 vccd1 vccd1 _11468_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12713__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13694__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ _06943_/A _13008_/X _13012_/X hold2774/X vssd1 vssd1 vccd1 vccd1 _13020_/A
+ sky130_fd_sc_hd__o211a_1
X_10225_ _10225_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10225_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10115__C _14959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10156_/A _10156_/B _10156_/C vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__or3_2
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14964_ _14971_/CLK _14964_/D vssd1 vssd1 vccd1 vccd1 _14964_/Q sky130_fd_sc_hd__dfxtp_2
X_10087_ _13885_/Q hold839/A hold685/A hold867/A _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _10087_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08089__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12572__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ _15448_/CLK _13915_/D vssd1 vssd1 vccd1 vccd1 _13915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10131__B _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14895_ _14989_/CLK _14895_/D vssd1 vssd1 vccd1 vccd1 _14895_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11942__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13846_ _14472_/CLK _13846_/D vssd1 vssd1 vccd1 vccd1 _13846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13442__B _13442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12720__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10989_ _10986_/X _10987_/Y _10805_/Y _10807_/X vssd1 vssd1 vccd1 vccd1 _10990_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12875__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12728_ _13519_/A0 _13103_/A2 _13078_/B1 _13188_/B vssd1 vssd1 vccd1 vccd1 _12728_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15447_ _15448_/CLK hold916/X vssd1 vssd1 vccd1 vccd1 hold915/A sky130_fd_sc_hd__dfxtp_1
X_12659_ hold1395/X hold2081/X _12866_/S vssd1 vssd1 vccd1 vccd1 _12659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12870__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15378_ _15378_/CLK hold378/X vssd1 vssd1 vccd1 vccd1 hold377/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14329_ _15292_/CLK _14329_/D vssd1 vssd1 vccd1 vccd1 _14329_/Q sky130_fd_sc_hd__dfxtp_1
Xhold405 hold405/A vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold416 hold416/A vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12074__A _14977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold438 hold438/A vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08702__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10306__B _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _09869_/A _09869_/B _09869_/C vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12802__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09383__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ _08820_/B _08820_/C _08820_/A vssd1 vssd1 vccd1 vccd1 _08821_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13617__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1105 _14744_/Q vssd1 vssd1 vccd1 vccd1 hold1105/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _07529_/X vssd1 vssd1 vccd1 vccd1 _14154_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ hold235/A _14311_/Q hold697/A _13971_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08752_/X sky130_fd_sc_hd__mux4_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 _14415_/Q vssd1 vssd1 vccd1 vccd1 hold1127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 _11937_/X vssd1 vssd1 vccd1 vccd1 _14757_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _14549_/Q vssd1 vssd1 vccd1 vccd1 hold1149/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__B2 _13178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07703_ hold627/X _11921_/A0 _07709_/S vssd1 vssd1 vccd1 vccd1 hold628/A sky130_fd_sc_hd__mux2_1
XANTENNA__07107__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08683_ _09661_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__and2_1
XFILLER_0_206_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11852__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07634_ hold1419/X _13740_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07634_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13417__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__S0 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _13396_/A hold181/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__and2_1
XANTENNA__09636__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A2 _13424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _09400_/B _09303_/C _09303_/A vssd1 vssd1 vccd1 vccd1 _09305_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11153__A _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07350__B _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__C1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ hold1169/X _13735_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07496_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ _14283_/Q _14219_/Q _14155_/Q hold873/A _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09236_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout607_A _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07777__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ _09016_/A _09015_/B _09013_/X vssd1 vssd1 vccd1 vccd1 _09178_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08117_ _08065_/A _08116_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08117_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12943__A1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08072__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__B _10010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _09514_/A _09096_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _09097_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_160_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__D _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08048_ _13546_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08257_/C sky130_fd_sc_hd__and2_1
XFILLER_0_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold950 hold950/A vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 hold961/A vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 hold972/A vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold983 hold983/A vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 hold994/A vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08375__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _10115_/B _10010_/B _10010_/C _10010_/D vssd1 vssd1 vccd1 vccd1 _10011_/B
+ sky130_fd_sc_hd__and4_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__C _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _11578_/A _10108_/C _14963_/Q _10000_/A vssd1 vssd1 vccd1 vccd1 _09999_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2340 hold2826/X vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__buf_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2351 hold2855/X vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__buf_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2362 _14974_/Q vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2373 _08004_/X vssd1 vssd1 vccd1 vccd1 hold2373/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2384 _14063_/Q vssd1 vssd1 vccd1 vccd1 _06922_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1650 _07699_/X vssd1 vssd1 vccd1 vccd1 _14319_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2395 _12195_/X vssd1 vssd1 vccd1 vccd1 _14908_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1661 _15427_/Q vssd1 vssd1 vccd1 vccd1 hold1661/X sky130_fd_sc_hd__dlygate4sd3_1
X_11961_ _13683_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__nor2_4
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09875__A1 _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1672 _07500_/X vssd1 vssd1 vccd1 vccd1 _14128_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1683 _14130_/Q vssd1 vssd1 vccd1 vccd1 hold1683/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1694 _07495_/X vssd1 vssd1 vccd1 vccd1 _14123_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11762__S _11762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _10910_/X _10912_/B vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__nand2b_1
X_13700_ hold405/X _13700_/A1 _13714_/S vssd1 vssd1 vccd1 vccd1 hold406/A sky130_fd_sc_hd__mux2_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _15454_/CLK _14680_/D vssd1 vssd1 vccd1 vccd1 _14680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ hold513/X _13746_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13631_ _09344_/A _13797_/A2 _13630_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _15343_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10843_ _11015_/B _10841_/Y _10619_/D _10620_/B vssd1 vssd1 vccd1 vccd1 _10844_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13562_ _14437_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13562_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12631__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ _11510_/A1 _10767_/Y _10769_/Y _10771_/Y _10773_/Y vssd1 vssd1 vccd1 vccd1
+ _10774_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08075__C _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13689__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15301_ _15301_/CLK _15301_/D vssd1 vssd1 vccd1 vccd1 _15301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ _12366_/A _12508_/X _12512_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12520_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _13495_/A hold133/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__and2_1
XFILLER_0_192_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_160_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15440_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08850__A2 _08851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07687__S _07693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _12644_/A1 _12439_/X _12443_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12445_/B
+ sky130_fd_sc_hd__o211a_1
X_15232_ _15243_/CLK _15232_/D vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _15426_/CLK _15163_/D vssd1 vssd1 vccd1 vccd1 _15163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12375_ _12692_/A1 _12372_/X _12374_/X vssd1 vssd1 vccd1 vccd1 _12375_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08602__A2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10945__B1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14114_ _15435_/CLK hold286/X vssd1 vssd1 vccd1 vccd1 _14114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ _11281_/A _11281_/B _11280_/A _11279_/Y vssd1 vssd1 vccd1 vccd1 _11471_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_120_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ _15383_/CLK hold394/X vssd1 vssd1 vccd1 vccd1 hold393/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10126__B _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12147__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__S _11943_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14045_ _14105_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11257_ _11254_/Y _11255_/X _11067_/X _11069_/Y vssd1 vssd1 vccd1 vccd1 _11258_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_24_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _10053_/Y _10055_/X _10206_/X _10207_/Y vssd1 vssd1 vccd1 vccd1 _10386_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13437__B _13437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _11614_/A _11542_/B _11564_/B _11586_/A vssd1 vssd1 vccd1 vccd1 _11188_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08461__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11238__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _10137_/X _10139_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10142__A _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13647__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__A1 _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14947_ _15293_/CLK _14947_/D vssd1 vssd1 vccd1 vccd1 _14947_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__08669__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14878_ _14992_/CLK _14878_/D vssd1 vssd1 vccd1 vccd1 _14878_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_187_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13172__B _13172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09618__A1 _11474_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ _15458_/CLK _13829_/D vssd1 vssd1 vccd1 vccd1 _13829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12848__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07350_ _10744_/A _15356_/Q _15340_/Q _15339_/Q vssd1 vssd1 vccd1 vccd1 _07351_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_0_70_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07281_ _08012_/B _10507_/A vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_151_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09020_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _09186_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07597__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09809__C _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2739_A _15180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__A2 _13398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09229__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13025__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11847__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13628__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09922_ _13750_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _09922_/Y sky130_fd_sc_hd__nor2_1
Xfanout704 _13691_/A1 vssd1 vssd1 vccd1 vccd1 _13724_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08357__A1 _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout715 hold479/X vssd1 vssd1 vccd1 vccd1 _13719_/A1 sky130_fd_sc_hd__buf_4
Xfanout726 _14960_/Q vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09853_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__nand2b_1
Xfanout737 _11390_/A vssd1 vssd1 vccd1 vccd1 _10316_/B sky130_fd_sc_hd__clkbuf_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _10306_/A vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__buf_4
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout759 _14949_/Q vssd1 vssd1 vccd1 vccd1 _11620_/A sky130_fd_sc_hd__clkbuf_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _08804_/A _08804_/B vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__xnor2_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _09918_/A _13446_/B _09783_/X vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__o21ai_1
X_06996_ _13668_/A1 hold1261/X _07010_/S vssd1 vssd1 vccd1 vccd1 _06996_/X sky130_fd_sc_hd__mux2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08735_ _11473_/A _08841_/B _08735_/C vssd1 vssd1 vccd1 vccd1 _08735_/X sky130_fd_sc_hd__and3_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09857__A1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13363__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _15209_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _08651_/Y _08656_/Y _08665_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08667_/B sky130_fd_sc_hd__a221o_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__B1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ hold913/X _13690_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 hold914/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08597_ _08597_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _08614_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_163_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout724_A _14962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07548_ _13386_/A hold211/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08293__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_142_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _14651_/CLK sky130_fd_sc_hd__clkbuf_16
X_07479_ hold895/X _13718_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 hold896/A sky130_fd_sc_hd__mux2_1
XFILLER_0_174_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12707__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _09218_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _13358_/B sky130_fd_sc_hd__nand2_1
X_10490_ _10652_/B _10489_/C _10489_/A vssd1 vssd1 vccd1 vccd1 _10491_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ _09033_/A _09032_/B _09032_/A vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08045__B1 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10927__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ _14891_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12160_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12129__C1 _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__S _11761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _11111_/A _11111_/B vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13538__A _15460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ hold2422/X _12099_/A2 _12090_/X _13495_/A vssd1 vssd1 vccd1 vccd1 _12091_/X
+ sky130_fd_sc_hd__o211a_1
Xhold780 hold780/A vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold791 hold791/A vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _11566_/A _15223_/Q _11229_/A _11042_/D vssd1 vssd1 vccd1 vccd1 _11229_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12775__S0 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07020__A1 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2170 _13521_/X vssd1 vssd1 vccd1 vccd1 _15279_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _15378_/CLK _14801_/D vssd1 vssd1 vccd1 vccd1 _14801_/Q sky130_fd_sc_hd__dfxtp_1
Xhold2181 _13924_/Q vssd1 vssd1 vccd1 vccd1 hold2181/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2192 _07461_/X vssd1 vssd1 vccd1 vccd1 _14091_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _13024_/S1 _12990_/X _12992_/X vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__a21o_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1480 _07146_/X vssd1 vssd1 vccd1 vccd1 _13956_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1491 _14553_/Q vssd1 vssd1 vccd1 vccd1 hold1491/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14732_ _15179_/CLK _14732_/D vssd1 vssd1 vccd1 vccd1 _14732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _13732_/A1 hold1799/X _11959_/S vssd1 vssd1 vccd1 vccd1 _11944_/X sky130_fd_sc_hd__mux2_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08367__A _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11875_ hold1915/X _13729_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11875_/X sky130_fd_sc_hd__mux2_1
X_14663_ _14775_/CLK hold966/X vssd1 vssd1 vccd1 vccd1 hold965/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _07430_/A _13625_/C _13613_/X _13622_/C1 vssd1 vssd1 vccd1 vccd1 _15334_/D
+ sky130_fd_sc_hd__o211a_1
X_10826_ _11542_/A _11536_/A _11588_/A _11623_/A vssd1 vssd1 vccd1 vccd1 _10826_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ _15042_/CLK _14594_/D vssd1 vssd1 vccd1 vccd1 _14594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10757_ hold157/A _14325_/Q hold623/A _13985_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10757_/X sky130_fd_sc_hd__mux4_1
X_13545_ _08038_/A _08441_/B _13544_/X _13178_/A vssd1 vssd1 vccd1 vccd1 _13545_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_133_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _15415_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13212__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _13481_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _15235_/D sky130_fd_sc_hd__and2_2
XFILLER_0_153_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10688_ _10688_/A _10688_/B vssd1 vssd1 vccd1 vccd1 _10691_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07210__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15215_ _15222_/CLK _15215_/D vssd1 vssd1 vccd1 vccd1 _15215_/Q sky130_fd_sc_hd__dfxtp_1
X_12427_ _13027_/A _12427_/B _12427_/C vssd1 vssd1 vccd1 vccd1 _12427_/X sky130_fd_sc_hd__and3_1
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput307 _14868_/Q vssd1 vssd1 vccd1 vccd1 out1[23] sky130_fd_sc_hd__buf_12
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _07907_/X _08636_/A _13141_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12359_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15146_ _15309_/CLK _15146_/D vssd1 vssd1 vccd1 vccd1 _15146_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput318 _14849_/Q vssd1 vssd1 vccd1 vccd1 out1[4] sky130_fd_sc_hd__buf_12
Xoutput329 _14827_/Q vssd1 vssd1 vccd1 vccd1 out2[14] sky130_fd_sc_hd__buf_12
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11667__S _11668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _11509_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15077_ _15077_/CLK hold528/X vssd1 vssd1 vccd1 vccd1 hold527/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ _13171_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _14938_/D sky130_fd_sc_hd__nor2_1
XANTENNA__07446__A _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ _14083_/CLK _14028_/D vssd1 vssd1 vccd1 vccd1 _14028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10697__A2 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11894__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__C _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08520_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08198__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13183__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09811__D _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2591_A _14993_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ _14791_/Q _14503_/Q _14631_/Q hold967/A _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08452_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_187_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07402_ _07402_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14032_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08382_ _08901_/A _08893_/A _09858_/A vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__and3_1
XFILLER_0_19_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07333_ _15338_/Q _15329_/Q _15328_/Q _15332_/Q vssd1 vssd1 vccd1 vccd1 _07334_/D
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13630__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15443_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12527__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07328_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09003_ _09571_/A _10126_/A _10126_/B _09435_/A vssd1 vssd1 vccd1 vccd1 _09003_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07120__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08027__B1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07195_ hold303/X _13663_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold304/A sky130_fd_sc_hd__mux2_1
XFILLER_0_131_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08578__A1 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13358__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _06943_/Y vssd1 vssd1 vccd1 vccd1 _13050_/S0 sky130_fd_sc_hd__buf_4
X_09905_ _09667_/Y _09670_/Y _09903_/A _09904_/X vssd1 vssd1 vccd1 vccd1 _09905_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 _10252_/A vssd1 vssd1 vccd1 vccd1 _08877_/A sky130_fd_sc_hd__clkbuf_4
Xfanout523 _08880_/A1 vssd1 vssd1 vccd1 vccd1 _06926_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout534 _15424_/Q vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__clkbuf_8
Xfanout545 _12211_/S1 vssd1 vssd1 vccd1 vccd1 _07815_/A sky130_fd_sc_hd__buf_4
Xfanout556 _15423_/Q vssd1 vssd1 vccd1 vccd1 _11501_/S1 sky130_fd_sc_hd__buf_4
X_09836_ _09833_/X _09834_/Y _09681_/B _09684_/B vssd1 vssd1 vccd1 vccd1 _09836_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout567 _10425_/S0 vssd1 vssd1 vccd1 vccd1 _10087_/S0 sky130_fd_sc_hd__buf_8
Xfanout578 _07448_/A vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__clkbuf_4
Xfanout589 _09809_/C vssd1 vssd1 vccd1 vccd1 _11378_/C sky130_fd_sc_hd__buf_6
XANTENNA__07790__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _09767_/A _09767_/B _09767_/C vssd1 vssd1 vccd1 vccd1 _09767_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_fanout841_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ _13651_/A1 hold1759/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06979_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11606__A _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08717_/B _08717_/C _08717_/A vssd1 vssd1 vccd1 vccd1 _08718_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _10000_/A _14961_/Q vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08649_ _13874_/Q hold303/A _13842_/Q _13810_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08649_/X sky130_fd_sc_hd__mux4_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _13691_/A1 hold1959/X _11668_/S vssd1 vssd1 vccd1 vccd1 _11660_/X sky130_fd_sc_hd__mux2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _10612_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10812_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11591_ _11589_/X _11441_/B _11591_/S vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_115_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15089_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11496__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13330_ input150/X fanout5/X fanout3/X input118/X vssd1 vssd1 vccd1 vccd1 _13330_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10542_ _10677_/A _10541_/C _10541_/A vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07030__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ input157/X fanout6/X fanout4/X input125/X vssd1 vssd1 vccd1 vccd1 _13261_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11060__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _11168_/A _11542_/A _11606_/A _11536_/A vssd1 vssd1 vccd1 vccd1 _10473_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_49_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13011__B1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12212_ _12247_/A _12212_/B vssd1 vssd1 vccd1 vccd1 _12212_/Y sky130_fd_sc_hd__nor2_1
X_15000_ _15254_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 _15000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12996__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _13396_/A _13192_/B vssd1 vssd1 vccd1 vccd1 _15057_/D sky130_fd_sc_hd__and2_1
XFILLER_0_60_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ hold2621/X _12173_/A2 _12142_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12143_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12748__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _14977_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12074_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_159_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10128__A1 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10404__B _10405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11025_ _11025_/A _11025_/B _11025_/C vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__and3_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10679__A2 _15219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13078__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__B _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13207__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10420__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _13101_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12977_/C sky130_fd_sc_hd__or2_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07205__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _15287_/CLK hold656/X vssd1 vssd1 vccd1 vccd1 hold655/A sky130_fd_sc_hd__dfxtp_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _13715_/A1 hold991/X _11927_/S vssd1 vssd1 vccd1 vccd1 hold992/A sky130_fd_sc_hd__mux2_1
XFILLER_0_185_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11950__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14646_ _15383_/CLK hold296/X vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11858_ hold651/X _13745_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold652/A sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13450__B _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _10806_/Y _10807_/X _10623_/C _10623_/Y vssd1 vssd1 vccd1 vccd1 _10810_/C
+ sky130_fd_sc_hd__o211ai_2
Xclkbuf_leaf_106_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _14989_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_19 _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ _15376_/CLK hold208/X vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11789_ hold485/X _11921_/A0 _11795_/S vssd1 vssd1 vccd1 vccd1 hold486/A sky130_fd_sc_hd__mux2_1
XANTENNA__08544__B _14434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _13742_/A1 hold2073/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_153_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13459_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _15223_/D sky130_fd_sc_hd__and2_1
XFILLER_0_152_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__A2 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_71_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13178__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15129_ _15132_/CLK _15129_/D vssd1 vssd1 vccd1 vccd1 _15129_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10017__D _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12739__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _07951_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07951_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10314__B _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_86_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _07882_/A _12252_/A _12252_/B vssd1 vssd1 vccd1 vccd1 _07882_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10033__C _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09621_ _11287_/S _09619_/Y _09767_/C _09618_/X vssd1 vssd1 vccd1 vccd1 _13393_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_128_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09552_ _09549_/X _09550_/Y _09408_/B _09411_/B vssd1 vssd1 vccd1 vccd1 _09552_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08503_ _08503_/A _08503_/B vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_195_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _12221_/B _09481_/Y _09619_/C _08526_/B hold2795/X vssd1 vssd1 vccd1 vccd1
+ _09483_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_188_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11860__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08434_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_144_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08735__A _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08365_ _08873_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _08365_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout422_A _13204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07316_ _15225_/Q _14969_/Q vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__or2_1
XFILLER_0_190_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ _08401_/B _08296_/B vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_117_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_159_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07247_ _10338_/C _11605_/B vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12691__S _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07785__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07178_ _13679_/A1 hold1403/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07178_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout791_A _13076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout889_A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08971__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__D _15354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout364 _12310_/X vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__buf_8
Xfanout375 _13502_/Y vssd1 vssd1 vccd1 vccd1 _13518_/S sky130_fd_sc_hd__clkbuf_16
Xfanout386 _11762_/S vssd1 vssd1 vccd1 vccd1 _11745_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_198_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09819_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__nor2_1
Xfanout397 _07610_/Y vssd1 vssd1 vccd1 vccd1 _07626_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12830_ _13080_/A1 _12829_/X _12827_/X vssd1 vssd1 vccd1 vccd1 _13160_/B sky130_fd_sc_hd__a21oi_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07025__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12917_/A1 _12760_/X _12844_/A1 vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12866__S _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14500_ _15365_/CLK _14500_/D vssd1 vssd1 vccd1 vccd1 _14500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11712_ hold669/X _13666_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold670/A sky130_fd_sc_hd__mux2_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12692_ _12692_/A1 _12691_/X _12366_/A vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__a21o_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11643_ _11643_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__nand2_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _15305_/CLK _14431_/D vssd1 vssd1 vccd1 vccd1 _14431_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11574_ _11574_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11575_/B sky130_fd_sc_hd__nand2_1
X_14362_ _15261_/CLK _14362_/D vssd1 vssd1 vccd1 vccd1 _14362_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10597__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 dmemresp_rdata[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
Xinput28 dmemresp_rdata[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13697__S _13698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13313_ input80/X fanout2/X _13312_/X vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__a21oi_1
Xinput39 imemresp_data[15] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
X_10525_ _11620_/A _11537_/B _10298_/X _10297_/X _11623_/A vssd1 vssd1 vccd1 vccd1
+ _10530_/A sky130_fd_sc_hd__a32o_1
X_14293_ _14776_/CLK _14293_/D vssd1 vssd1 vccd1 vccd1 _14293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07695__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13244_ input65/X fanout1/X _13243_/X vssd1 vssd1 vccd1 vccd1 _13245_/B sky130_fd_sc_hd__a21oi_1
X_10456_ _11590_/A _11573_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _10456_/X sky130_fd_sc_hd__and3_1
XANTENNA_output174_A _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07214__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13175_ _13477_/A _13175_/B vssd1 vssd1 vccd1 vccd1 _15040_/D sky130_fd_sc_hd__and2_1
XFILLER_0_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _10387_/A _10387_/B _10387_/C vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _15003_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12126_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10134__B _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _12059_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _14841_/D sky130_fd_sc_hd__and2_1
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ _11564_/A _11378_/C _11010_/C _11010_/D vssd1 vssd1 vccd1 vccd1 _11008_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07443__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08478__B1 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12959_ hold833/X hold2211/X _13066_/S vssd1 vssd1 vccd1 vccd1 _12959_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11680__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08555__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13180__B _13180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14629_ _14783_/CLK hold376/X vssd1 vssd1 vccd1 vccd1 hold375/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09978__B1 _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _08149_/B _08149_/C _08149_/A vssd1 vssd1 vccd1 vccd1 _08152_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11412__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07101_ _13737_/A1 hold1875/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07101_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08876__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08081_ _08080_/A _08080_/B _08080_/C vssd1 vssd1 vccd1 vccd1 _08082_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08650__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09386__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07032_ hold565/X _13703_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold566/A sky130_fd_sc_hd__mux2_1
XFILLER_0_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08290__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _12241_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08983_/Y sky130_fd_sc_hd__nor2_1
Xhold2703 _15183_/Q vssd1 vssd1 vccd1 vccd1 hold2703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2714 _15129_/Q vssd1 vssd1 vccd1 vccd1 _06941_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10760__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2725 _12026_/X vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13636__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2736 _15123_/Q vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__dlygate4sd3_1
X_07934_ _08197_/A _07934_/B vssd1 vssd1 vccd1 vccd1 _07934_/X sky130_fd_sc_hd__or2_1
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2747 _15181_/Q vssd1 vssd1 vccd1 vccd1 hold2747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2758 _15106_/Q vssd1 vssd1 vccd1 vccd1 hold2758/X sky130_fd_sc_hd__buf_1
XFILLER_0_208_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2769 _15196_/Q vssd1 vssd1 vccd1 vccd1 hold2769/X sky130_fd_sc_hd__buf_1
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07865_ _07863_/Y _07864_/X _14093_/Q _06972_/B vssd1 vssd1 vccd1 vccd1 _07865_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10512__A1 _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout372_A _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__C _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _09461_/C _09464_/B _09601_/X _09603_/Y vssd1 vssd1 vccd1 vccd1 _09604_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_78_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07796_ hold977/X _13734_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold978/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09535_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout637_A _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10276__B1 _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09317_/X _09321_/B _09463_/X _09465_/Y vssd1 vssd1 vccd1 vccd1 _09466_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__12360__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07141__A0 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08417_ _08322_/A _08322_/C _08322_/B vssd1 vssd1 vccd1 vccd1 _08418_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _10351_/A _11536_/B _09398_/A vssd1 vssd1 vccd1 vccd1 _09397_/X sky130_fd_sc_hd__and3_1
XFILLER_0_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout804_A _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08348_ _15141_/Q _11643_/B _07390_/A vssd1 vssd1 vccd1 vccd1 _08348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10579__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08867__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08279_ _14661_/Q _13934_/Q _15435_/Q _13902_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08280_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10310_ _10308_/X _10310_/B vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ _11645_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11290_/Y sky130_fd_sc_hd__nor2_1
X_10241_ _10244_/A _10238_/X _10240_/X vssd1 vssd1 vccd1 vccd1 _10241_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10172_ _10172_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11765__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14980_ _15248_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 _14980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13931_ _15432_/CLK _13931_/D vssd1 vssd1 vccd1 vccd1 _13931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__B _14971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13862_ _15296_/CLK _13862_/D vssd1 vssd1 vccd1 vccd1 _13862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__A2 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ _12917_/B1 _12808_/X _12812_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12820_/A
+ sky130_fd_sc_hd__o211a_1
X_13793_ hold2569/X _13797_/A2 _13626_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15422_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13281__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10806__A2 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12744_ _12844_/A1 hold2806/X _12743_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12744_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12671_/X _12672_/X _12674_/X _12673_/X _12700_/S0 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12676_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_167_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14414_ _15410_/CLK hold644/X vssd1 vssd1 vccd1 vccd1 hold643/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11626_ _11626_/A _11626_/B _11626_/C vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__and3_1
XFILLER_0_182_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15394_ _15394_/CLK _15394_/D vssd1 vssd1 vccd1 vccd1 _15394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10129__B _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14345_ _14409_/CLK hold464/X vssd1 vssd1 vccd1 vccd1 hold463/A sky130_fd_sc_hd__dfxtp_1
X_11557_ _11557_/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09918__B _13448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13220__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10508_ _11550_/A _11614_/B _11586_/B _10507_/A vssd1 vssd1 vccd1 vccd1 _10510_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 hold609/A vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
X_11488_ hold2328/X _07812_/A _13636_/B _11485_/Y _11487_/X vssd1 vssd1 vccd1 vccd1
+ _11488_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14276_ _15437_/CLK hold822/X vssd1 vssd1 vccd1 vccd1 hold821/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10439_ _10439_/A _10439_/B vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__nor2_1
X_13227_ hold837/X _13673_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold838/A sky130_fd_sc_hd__mux2_1
XFILLER_0_21_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09934__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12731__A2 _13156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _13389_/A _13158_/B vssd1 vssd1 vccd1 vccd1 _15023_/D sky130_fd_sc_hd__nor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11675__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ hold2455/X _12129_/A2 _12108_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12109_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13456__A _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13089_ _14297_/Q _14233_/Q _14169_/Q _14487_/Q _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13089_/X sky130_fd_sc_hd__mux4_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1309 _14752_/Q vssd1 vssd1 vccd1 vccd1 hold1309/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10799__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09360__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07650_ hold503/X _13689_/A1 _07660_/S vssd1 vssd1 vccd1 vccd1 hold504/A sky130_fd_sc_hd__mux2_1
XFILLER_0_178_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11407__C _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07581_ _13687_/A1 hold1739/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09320_ _09316_/Y _09318_/X _09184_/B _09186_/B vssd1 vssd1 vccd1 vccd1 _09321_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__09112__A1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13191__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08285__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _09435_/A _09864_/C _09714_/D _09253_/A vssd1 vssd1 vccd1 vccd1 _09255_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07674__A1 _15066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold2769_A _15196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ hold519/A hold901/A hold543/A _14756_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08202_/X sky130_fd_sc_hd__mux4_1
X_09182_ _09049_/X _09051_/Y _09180_/X _09181_/Y vssd1 vssd1 vccd1 vccd1 _09184_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11758__A0 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08133_ _08118_/Y _08123_/Y _08132_/X _08760_/A _12252_/A vssd1 vssd1 vccd1 vccd1
+ _08134_/B sky130_fd_sc_hd__a221o_1
XANTENNA__09828__B _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_6__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_08064_ hold435/A _13931_/Q hold661/A _13899_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08065_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10430__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10981__A1 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07015_ hold859/X _13719_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 hold860/A sky130_fd_sc_hd__mux2_1
XFILLER_0_141_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07348__B _15354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout587_A _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2500 _10413_/X vssd1 vssd1 vccd1 vccd1 _14448_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13366__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2511 _14846_/Q vssd1 vssd1 vccd1 vccd1 hold2511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2522 _12268_/B vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2533 _08645_/Y vssd1 vssd1 vccd1 vccd1 hold2533/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12270__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _08966_/A _09346_/B _08966_/C vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__or3_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2544 hold2829/X vssd1 vssd1 vccd1 vccd1 _11291_/B sky130_fd_sc_hd__clkbuf_2
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1810 _11823_/X vssd1 vssd1 vccd1 vccd1 _14647_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2555 _14998_/Q vssd1 vssd1 vccd1 vccd1 hold2555/X sky130_fd_sc_hd__buf_2
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2566 _15355_/Q vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__clkbuf_4
X_07917_ _06905_/A _07431_/A _08036_/S vssd1 vssd1 vccd1 vccd1 _07919_/B sky130_fd_sc_hd__mux2_2
Xhold1821 _14282_/Q vssd1 vssd1 vccd1 vccd1 hold1821/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12486__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1832 _07614_/X vssd1 vssd1 vccd1 vccd1 _14237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2577 _11118_/X vssd1 vssd1 vccd1 vccd1 _14452_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2588 _15111_/Q vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08897_ _08780_/X _08782_/X _08895_/Y _08896_/X vssd1 vssd1 vccd1 vccd1 _08897_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout754_A _14950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1843 _15403_/Q vssd1 vssd1 vccd1 vccd1 hold1843/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08154__A2 _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1854 _07197_/X vssd1 vssd1 vccd1 vccd1 _14004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_95_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15251_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2599 _07982_/X vssd1 vssd1 vccd1 vccd1 _14427_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1865 _14406_/Q vssd1 vssd1 vccd1 vccd1 hold1865/X sky130_fd_sc_hd__dlygate4sd3_1
X_07848_ hold195/A hold95/A hold197/A _07847_/X _14057_/Q vssd1 vssd1 vccd1 vccd1
+ _07848_/X sky130_fd_sc_hd__o41a_1
Xhold1876 _07101_/X vssd1 vssd1 vccd1 vccd1 _13914_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1887 _13996_/Q vssd1 vssd1 vccd1 vccd1 hold1887/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1898 _11921_/X vssd1 vssd1 vccd1 vccd1 _14742_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10592__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__A2 _13376_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__A1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07779_ hold591/X _12329_/A _07794_/S vssd1 vssd1 vccd1 vccd1 hold592/A sky130_fd_sc_hd__mux2_1
XFILLER_0_196_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11614__A _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09518_ _09503_/Y _09508_/Y _09517_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09519_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ _10790_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10792_/B sky130_fd_sc_hd__xor2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08195__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09654__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11333__B _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A _09449_/B _09449_/C vssd1 vssd1 vccd1 vccd1 _09450_/B sky130_fd_sc_hd__nor3_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _14659_/Q _13932_/Q _12460_/S vssd1 vssd1 vccd1 vccd1 _12460_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11749__A0 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11411_ _11563_/A _11569_/B _11563_/B _11594_/A vssd1 vssd1 vccd1 vccd1 _11414_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12391_ hold595/A _14237_/Q _12460_/S vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13040__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11342_ _11343_/A _11343_/B _11343_/C vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__o21a_1
X_14130_ _15093_/CLK _14130_/D vssd1 vssd1 vccd1 vccd1 _14130_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08090__A1 _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11273_ _11273_/A _11273_/B _11273_/C vssd1 vssd1 vccd1 vccd1 _11273_/Y sky130_fd_sc_hd__nor3_1
X_14061_ _15348_/CLK _14061_/D vssd1 vssd1 vccd1 vccd1 _14061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10224_ _07320_/D _07302_/B _10077_/B _11640_/B1 vssd1 vssd1 vccd1 vccd1 _10225_/B
+ sky130_fd_sc_hd__a31o_1
X_13012_ _13099_/S1 _13009_/X _13011_/X vssd1 vssd1 vccd1 vccd1 _13012_/X sky130_fd_sc_hd__a21o_1
X_10155_ _10154_/B _10154_/C _10154_/A vssd1 vssd1 vccd1 vccd1 _10156_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__10115__D _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ _14971_/CLK _14963_/D vssd1 vssd1 vccd1 vccd1 _14963_/Q sky130_fd_sc_hd__dfxtp_4
X_10086_ hold269/A hold335/A _14612_/Q _13981_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _10086_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08089__B _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15246_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09342__A1 _11287_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ _15411_/CLK _13914_/D vssd1 vssd1 vccd1 vccd1 _13914_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12572__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__C _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14894_ _14989_/CLK _14894_/D vssd1 vssd1 vccd1 vccd1 _14894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13845_ _14602_/CLK _13845_/D vssd1 vssd1 vccd1 vccd1 _13845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13215__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ hold207/X vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__clkbuf_1
X_10988_ _10805_/Y _10807_/X _10986_/X _10987_/Y vssd1 vssd1 vccd1 vccd1 _10990_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07213__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _13102_/A _12727_/B _12727_/C vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__and3_1
XFILLER_0_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15446_ _15446_/CLK hold512/X vssd1 vssd1 vccd1 vccd1 hold511/A sky130_fd_sc_hd__dfxtp_1
X_12658_ hold909/X hold653/X hold1015/X hold1297/X _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12658_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12456__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ _11609_/A _11609_/B vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__xor2_1
X_15377_ _15377_/CLK hold696/X vssd1 vssd1 vccd1 vccd1 hold695/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12589_ hold993/A _14213_/Q _14149_/Q _14467_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12589_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15315_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _14651_/CLK _14328_/D vssd1 vssd1 vccd1 vccd1 _14328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold406 hold406/A vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 hold417/A vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold428 hold428/A vssd1 vssd1 vccd1 vccd1 hold428/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold439 hold439/A vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14259_ _14419_/CLK hold568/X vssd1 vssd1 vccd1 vccd1 hold567/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07883__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12704__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ _08820_/A _08820_/B _08820_/C vssd1 vssd1 vccd1 vccd1 _08820_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__13186__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__B _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__A _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_99_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _11923_/X vssd1 vssd1 vccd1 vccd1 _14744_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _14730_/Q vssd1 vssd1 vccd1 vccd1 hold1117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 _07800_/X vssd1 vssd1 vccd1 vccd1 _14415_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ _13570_/B _08749_/Y _08750_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _08751_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 _13858_/Q vssd1 vssd1 vccd1 vccd1 hold1139/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_77_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15458_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08136__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08767__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ hold297/X _13675_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08682_ _09816_/A _09858_/C vssd1 vssd1 vccd1 vccd1 _08692_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__B2 _13201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07633_ hold699/X _13739_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold700/A sky130_fd_sc_hd__mux2_1
XANTENNA__12545__C_N _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07564_ _13396_/A hold139/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__and2_1
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12315__S1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07123__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09303_ _09303_/A _09400_/B _09303_/C vssd1 vssd1 vccd1 vccd1 _09305_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11153__B _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ hold1693/X _13734_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07495_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12581__A1_N _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12695__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _09941_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ _09165_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09078__A1_N _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout502_A _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12265__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ _13868_/Q _13996_/Q _13836_/Q _13804_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08116_/X sky130_fd_sc_hd__mux4_1
X_09096_ _13878_/Q _14006_/Q _13846_/Q _13814_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09096_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08072__B2 _13177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08047_ _14428_/Q _08441_/B _08034_/Y _08046_/X _13178_/A vssd1 vssd1 vccd1 vccd1
+ _08047_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_101_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold940 hold940/A vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 hold951/A vssd1 vssd1 vccd1 vccd1 hold951/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07793__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold962 hold962/A vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 hold973/A vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 hold984/A vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 hold995/A vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12204__S _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ _09997_/B _09997_/C _09997_/A vssd1 vssd1 vccd1 vccd1 _10056_/B sky130_fd_sc_hd__a21o_1
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__D _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2330 _11489_/X vssd1 vssd1 vccd1 vccd1 _14454_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2341 _14029_/Q vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2352 _14991_/Q vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__buf_2
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _08948_/B _08948_/C _08948_/A vssd1 vssd1 vccd1 vccd1 _08950_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2363 _12135_/X vssd1 vssd1 vccd1 vccd1 _14878_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _14909_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2374 _08033_/Y vssd1 vssd1 vccd1 vccd1 _13414_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1640 _07174_/X vssd1 vssd1 vccd1 vccd1 _13982_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2385 _14429_/Q vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_93_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1651 _14504_/Q vssd1 vssd1 vccd1 vccd1 hold1651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2396 hold2847/X vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__buf_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1662 _13717_/X vssd1 vssd1 vccd1 vccd1 _15427_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ _13715_/A1 hold1389/X _11960_/S vssd1 vssd1 vccd1 vccd1 _11960_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_169_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1673 _14679_/Q vssd1 vssd1 vccd1 vccd1 hold1673/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08918__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__A2 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1684 _07502_/X vssd1 vssd1 vccd1 vccd1 _14130_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _10726_/Y _10730_/A _11098_/B _10909_/X vssd1 vssd1 vccd1 vccd1 _10912_/B
+ sky130_fd_sc_hd__a211o_1
Xhold1695 _14207_/Q vssd1 vssd1 vccd1 vccd1 hold1695/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ hold731/X _13745_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 hold732/A sky130_fd_sc_hd__mux2_1
XANTENNA__13035__S _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ input41/X _13634_/B vssd1 vssd1 vccd1 vccd1 _13630_/X sky130_fd_sc_hd__or2_1
X_10842_ _10619_/D _10620_/B _11015_/B _10841_/Y vssd1 vssd1 vccd1 vccd1 _10844_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07033__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12631__A1 _13106_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _08743_/A _09222_/B _13560_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _13561_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10773_ _11493_/A _10772_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _10773_/Y sky130_fd_sc_hd__o21ai_1
X_15300_ _15301_/CLK _15300_/D vssd1 vssd1 vccd1 vccd1 _15300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08075__D _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__S _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _12368_/A _12509_/X _12511_/X vssd1 vssd1 vccd1 vccd1 _12512_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_164_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _13492_/A hold57/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__and2_1
XFILLER_0_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12919__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15231_ _15251_/CLK _15231_/D vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
X_12443_ _12474_/S1 _12440_/X _12442_/X vssd1 vssd1 vccd1 vccd1 _12443_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07269__A _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15162_ _15296_/CLK _15162_/D vssd1 vssd1 vccd1 vccd1 _15162_/Q sky130_fd_sc_hd__dfxtp_1
X_12374_ _12668_/A1 _12373_/X _12366_/A vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ _15040_/CLK _14113_/D vssd1 vssd1 vccd1 vccd1 _14113_/Q sky130_fd_sc_hd__dfxtp_1
X_11325_ _07240_/B _07328_/A _11323_/X _11640_/B1 vssd1 vssd1 vccd1 vccd1 _11325_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15093_ _15093_/CLK hold742/X vssd1 vssd1 vccd1 vccd1 hold741/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__C _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14044_ _14105_/CLK hold198/X vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__dfxtp_1
X_11256_ _11067_/X _11069_/Y _11254_/Y _11255_/X vssd1 vssd1 vccd1 vccd1 _11329_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12242__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output254_A _14428_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09563__A1 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10207_ _10206_/A _10206_/B _10206_/C _10206_/D vssd1 vssd1 vccd1 vccd1 _10207_/Y
+ sky130_fd_sc_hd__o22ai_2
X_11187_ _11183_/Y _11184_/X _10996_/A _10996_/Y vssd1 vssd1 vccd1 vccd1 _11220_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07208__S _07214_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10138_ _10135_/Y _10136_/X _10024_/C _10023_/Y vssd1 vssd1 vccd1 vccd1 _10139_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11238__B _15226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__B _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15132_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11953__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10069_ _10266_/B _10263_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__or2_1
X_14946_ _15225_/CLK _14946_/D vssd1 vssd1 vccd1 vccd1 _14946_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11122__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14877_ _15248_/CLK _14877_/D vssd1 vssd1 vccd1 vccd1 _14877_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13828_ _15384_/CLK _13828_/D vssd1 vssd1 vccd1 vccd1 _13828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07629__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ hold203/X vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__12784__S _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07280_ _07280_/A _07280_/B vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15429_ _15429_/CLK hold636/X vssd1 vssd1 vccd1 vccd1 hold635/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12386__B1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__D _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08054__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10936__A1 _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09229__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _09929_/B _09921_/B vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09003__B1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13628__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout705 _15044_/Q vssd1 vssd1 vccd1 vccd1 _13691_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11429__A _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__S0 _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 _13652_/A1 vssd1 vssd1 vccd1 vccd1 _13718_/A1 sky130_fd_sc_hd__buf_4
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout727 _14960_/Q vssd1 vssd1 vccd1 vccd1 _10115_/D sky130_fd_sc_hd__buf_4
XANTENNA__12333__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 _14955_/Q vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__clkbuf_8
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 _10306_/A vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__clkbuf_4
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07118__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ _09164_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _13750_/A _13362_/B _09781_/X _09782_/Y vssd1 vssd1 vccd1 vccd1 _09783_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12959__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06995_ _13519_/A0 hold1035/X _07010_/S vssd1 vssd1 vccd1 vccd1 _06995_/X sky130_fd_sc_hd__mux2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11863__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _08734_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _08735_/C sky130_fd_sc_hd__or2_1
XANTENNA__09857__A2 _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _08992_/A1 _08658_/Y _08660_/Y _08662_/Y _08664_/Y vssd1 vssd1 vccd1 vccd1
+ _08665_/X sky130_fd_sc_hd__o32a_1
XANTENNA__12861__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_109 _15209_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07616_ hold1991/X _13689_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07616_/X sky130_fd_sc_hd__mux2_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _10351_/A _09858_/C _08597_/A vssd1 vssd1 vccd1 vccd1 _08596_/X sky130_fd_sc_hd__and3_1
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07547_ _13386_/A hold189/X vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__and2_1
XANTENNA__12613__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07788__S _07794_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08293__A1 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ hold985/X _12329_/A _07493_/S vssd1 vssd1 vccd1 vccd1 hold986/A sky130_fd_sc_hd__mux2_1
XANTENNA__08293__B2 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _09217_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__or2_1
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08045__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _09317_/A _09148_/B vssd1 vssd1 vccd1 vccd1 _09190_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12472__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09793__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _13389_/B vssd1 vssd1 vccd1 vccd1 _09079_/Y sky130_fd_sc_hd__inv_2
X_11110_ _11110_/A _11110_/B vssd1 vssd1 vccd1 vccd1 _11111_/B sky130_fd_sc_hd__nor2_1
X_12090_ _14985_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12090_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__07817__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13538__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 hold770/A vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 hold781/A vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _11333_/B _15221_/Q _15222_/Q _11526_/A vssd1 vssd1 vccd1 vccd1 _11042_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08348__A2 _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold792 hold792/A vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12775__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07028__S _07028_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2160 _11954_/X vssd1 vssd1 vccd1 vccd1 _14774_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11773__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _15056_/CLK hold456/X vssd1 vssd1 vccd1 vccd1 hold455/A sky130_fd_sc_hd__dfxtp_1
Xhold2171 _14479_/Q vssd1 vssd1 vccd1 vccd1 hold2171/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2182 _07111_/X vssd1 vssd1 vccd1 vccd1 _13924_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2193 _13824_/Q vssd1 vssd1 vccd1 vccd1 hold2193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12992_ _13092_/A1 _12991_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _12992_/X sky130_fd_sc_hd__a21o_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07552__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 _13708_/X vssd1 vssd1 vccd1 vccd1 _15414_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1481 _13822_/Q vssd1 vssd1 vccd1 vccd1 hold1481/X sky130_fd_sc_hd__dlygate4sd3_1
X_14731_ _14731_/CLK _14731_/D vssd1 vssd1 vccd1 vccd1 _14731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1492 _11759_/X vssd1 vssd1 vccd1 vccd1 _14553_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11943_ _13698_/A1 hold1297/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14662_ _15436_/CLK _14662_/D vssd1 vssd1 vccd1 vccd1 _14662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11874_ hold1385/X _13728_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ input63/X _13636_/B vssd1 vssd1 vccd1 vccd1 _13613_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08808__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _10825_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _10835_/A sky130_fd_sc_hd__xor2_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12604__A1 _13385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14593_ _14595_/CLK hold862/X vssd1 vssd1 vccd1 vccd1 hold861/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07698__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ _14428_/Q _13554_/B vssd1 vssd1 vccd1 vccd1 _13544_/X sky130_fd_sc_hd__or2_1
XANTENNA__08383__A _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__B2 _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _13588_/A _13591_/A2 _10755_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _10756_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13475_ _13481_/A _13475_/B vssd1 vssd1 vccd1 vccd1 _13475_/X sky130_fd_sc_hd__and2_1
X_10687_ _11340_/A _15222_/Q vssd1 vssd1 vccd1 vccd1 _10688_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15214_ _15214_/CLK _15214_/D vssd1 vssd1 vccd1 vccd1 _15214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13565__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ _12676_/A _12426_/B vssd1 vssd1 vccd1 vccd1 _12427_/C sky130_fd_sc_hd__or2_1
XFILLER_0_23_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11948__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput308 _14869_/Q vssd1 vssd1 vccd1 vccd1 out1[24] sky130_fd_sc_hd__buf_12
X_15145_ _15309_/CLK _15145_/D vssd1 vssd1 vccd1 vccd1 _15145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _13027_/A _12353_/X _12356_/X vssd1 vssd1 vccd1 vccd1 _13141_/B sky130_fd_sc_hd__a21oi_4
Xoutput319 _14850_/Q vssd1 vssd1 vccd1 vccd1 out1[5] sky130_fd_sc_hd__buf_12
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _11497_/A _11305_/X _11307_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _11309_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13448__B _13448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15076_ _15365_/CLK _15076_/D vssd1 vssd1 vccd1 vccd1 _15076_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12215__S0 _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12288_ _13479_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _14937_/D sky130_fd_sc_hd__and2_1
X_14027_ _14083_/CLK hold256/X vssd1 vssd1 vccd1 vccd1 _14027_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07446__B _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _11239_/A _11239_/B vssd1 vssd1 vccd1 vccd1 _11258_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11683__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__D _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13464__A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__B _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08198__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14929_ _15243_/CLK _14929_/D vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12843__A1 _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08450_ _15368_/Q _15271_/Q _15079_/Q _14372_/Q _07816_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08450_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07401_ _07401_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14031_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08381_ _08893_/A _09860_/A _09858_/A _08901_/A vssd1 vssd1 vccd1 vccd1 _08384_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07332_ _13535_/A _07332_/B _12221_/A vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__and3_4
XFILLER_0_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ _15227_/Q _14971_/Q vssd1 vssd1 vccd1 vccd1 _07264_/B sky130_fd_sc_hd__or2_1
XFILLER_0_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ _09714_/A _10129_/A vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07194_ hold891/X _13662_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold892/A sky130_fd_sc_hd__mux2_1
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11858__S _11861_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08740__B _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12262__B _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ _09900_/Y _09901_/X _09747_/X _09749_/Y vssd1 vssd1 vccd1 vccd1 _09904_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout502 _12692_/A1 vssd1 vssd1 vccd1 vccd1 _12642_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout513 _09514_/A vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__buf_6
Xfanout524 _15425_/Q vssd1 vssd1 vccd1 vccd1 _08880_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12531__B1 _13148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 _15424_/Q vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__buf_6
XANTENNA__10768__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 _15423_/Q vssd1 vssd1 vccd1 vccd1 _12211_/S1 sky130_fd_sc_hd__clkbuf_4
X_09835_ _09681_/B _09684_/B _09833_/X _09834_/Y vssd1 vssd1 vccd1 vccd1 _09835_/Y
+ sky130_fd_sc_hd__a211oi_4
Xfanout557 _08763_/S0 vssd1 vssd1 vccd1 vccd1 _08548_/S0 sky130_fd_sc_hd__buf_8
Xfanout568 _10425_/S0 vssd1 vssd1 vccd1 vccd1 _09795_/S0 sky130_fd_sc_hd__buf_8
Xfanout579 _15220_/Q vssd1 vssd1 vccd1 vccd1 _11620_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout667_A _15062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13374__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09766_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13087__A1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ _07182_/A _11928_/A vssd1 vssd1 vccd1 vccd1 _06978_/X sky130_fd_sc_hd__or2_4
X_08717_ _08717_/A _08717_/B _08717_/C vssd1 vssd1 vccd1 vccd1 _08717_/Y sky130_fd_sc_hd__nand3_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__B _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09697_ _09693_/A _09694_/Y _09555_/B _09557_/B vssd1 vssd1 vccd1 vccd1 _09745_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout834_A _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ hold247/A hold365/A _14601_/Q _13970_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08648_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10940__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _08709_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _08617_/A sky130_fd_sc_hd__or2_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _11577_/A _11594_/B _10440_/X _10273_/B _14966_/Q vssd1 vssd1 vccd1 vccd1
+ _10612_/B sky130_fd_sc_hd__a32o_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11590_ _11590_/A _14966_/Q vssd1 vssd1 vccd1 vccd1 _11591_/S sky130_fd_sc_hd__nand2_1
XANTENNA__11496__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10541_ _10541_/A _10677_/A _10541_/C vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13547__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ _13287_/A _13260_/B vssd1 vssd1 vccd1 vccd1 _15106_/D sky130_fd_sc_hd__nor2_1
XANTENNA__11060__C _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13011__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10472_ _10472_/A _10472_/B vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_134_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11768__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ hold619/A _14202_/Q hold391/A _14456_/Q _12198_/S _12211_/S1 vssd1 vssd1
+ vccd1 vccd1 _12212_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_161_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _13397_/A _13191_/B vssd1 vssd1 vccd1 vccd1 _15056_/D sky130_fd_sc_hd__and2_1
XANTENNA__12996__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08974__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _14882_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12142_/X sky130_fd_sc_hd__or2_1
XFILLER_0_209_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09518__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12748__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ hold2513/X _12099_/A2 _12072_/X _13492_/A vssd1 vssd1 vccd1 vccd1 _12073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09762__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ _10844_/A _10844_/C _10844_/B vssd1 vssd1 vccd1 vccd1 _11025_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13284__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13078__B2 _13202_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__A _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12971_/X _12972_/X _12974_/X _12973_/X _13100_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _12976_/B sky130_fd_sc_hd__mux4_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _15418_/CLK hold514/X vssd1 vssd1 vccd1 vccd1 hold513/A sky130_fd_sc_hd__dfxtp_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _13681_/A1 hold2269/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _15093_/CLK hold920/X vssd1 vssd1 vccd1 vccd1 hold919/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ hold1773/X _13744_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 _11857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13223__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _10623_/C _10623_/Y _10806_/Y _10807_/X vssd1 vssd1 vccd1 vccd1 _10978_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13250__A1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14576_ _15444_/CLK hold218/X vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__dfxtp_1
X_11788_ hold311/X _13675_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold312/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13527_ _13675_/A1 hold625/X _13534_/S vssd1 vssd1 vccd1 vccd1 hold626/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10739_ _10958_/A _10737_/X _10738_/Y vssd1 vssd1 vccd1 vccd1 _10739_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13458_ _10744_/B _12286_/B _13466_/A vssd1 vssd1 vccd1 vccd1 _13459_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_152_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11678__S _11684_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ hold811/X hold1563/X _12459_/S vssd1 vssd1 vccd1 vccd1 _12409_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13553__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13459__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13389_ _13389_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _15180_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12761__B1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15128_ _15132_/CLK _15128_/D vssd1 vssd1 vccd1 vccd1 _15128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13178__B _13178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07950_ _07237_/B _07887_/B _08007_/A vssd1 vssd1 vccd1 vccd1 _07951_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12739__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15059_ _15449_/CLK _15059_/D vssd1 vssd1 vccd1 vccd1 _15059_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10314__C _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07881_ _07899_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__nand2b_4
XANTENNA__10033__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _09619_/B _09619_/C _09619_/A vssd1 vssd1 vccd1 vccd1 _09767_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13194__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__A1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _09408_/B _09411_/B _09549_/X _09550_/Y vssd1 vssd1 vccd1 vccd1 _09551_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08502_ _08502_/A _08502_/B vssd1 vssd1 vccd1 vccd1 _08598_/B sky130_fd_sc_hd__or2_1
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09482_ _07243_/B _09340_/A _09340_/B _09481_/A _07241_/Y vssd1 vssd1 vccd1 vccd1
+ _09619_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _08347_/A _08344_/Y _08346_/B vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08364_ hold499/A _14243_/Q hold925/A _14115_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08365_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12675__S0 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07131__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07315_ _07313_/X _08338_/C vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13792__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08295_ _08776_/A _08926_/A _08294_/C _08294_/D vssd1 vssd1 vccd1 vccd1 _08296_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout415_A _13716_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07246_ _09133_/A _08528_/D vssd1 vssd1 vccd1 vccd1 _08340_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13369__A _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ _13744_/A1 hold1177/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07177_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12201__C1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12273__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout784_A _14942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08971__A2 _13434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09582__A _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout365 _07903_/Y vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__buf_4
Xfanout376 _13502_/Y vssd1 vssd1 vccd1 vccd1 _13534_/S sky130_fd_sc_hd__clkbuf_16
X_09818_ _09666_/A _09665_/B _09665_/A vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout387 _11696_/Y vssd1 vssd1 vccd1 vccd1 _11712_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__10521__A _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _07610_/Y vssd1 vssd1 vccd1 vccd1 _07642_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_0_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09359__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _09557_/X _09602_/A _09747_/X _09748_/Y vssd1 vssd1 vccd1 vccd1 _09749_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12760_ _14671_/Q _13944_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__mux2_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__A _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07830__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ hold1205/X _13665_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ hold463/A hold601/A _12741_/S vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_210_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11352__A _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14430_ _15305_/CLK _14430_/D vssd1 vssd1 vccd1 vccd1 _14430_/Q sky130_fd_sc_hd__dfxtp_2
X_11642_ _07879_/X _11641_/X _11514_/X vssd1 vssd1 vccd1 vccd1 _13468_/B sky130_fd_sc_hd__a21oi_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13232__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07041__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14361_ _15292_/CLK _14361_/D vssd1 vssd1 vccd1 vccd1 _14361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput18 dmemresp_rdata[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
X_13312_ input144/X fanout5/X fanout3/X input112/X vssd1 vssd1 vccd1 vccd1 _13312_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10532_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 dmemresp_rdata[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_2
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14292_ _14775_/CLK _14292_/D vssd1 vssd1 vccd1 vccd1 _14292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13243_ input129/X fanout6/X fanout4/X input97/X vssd1 vssd1 vccd1 vccd1 _13243_/X
+ sky130_fd_sc_hd__a22o_1
X_10455_ _10455_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_33_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13174_ _13481_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _15039_/D sky130_fd_sc_hd__and2_1
X_10386_ _10386_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10387_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_21_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output167_A _15179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__A2 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ hold2518/X _12129_/A2 _12124_/X _12063_/A vssd1 vssd1 vccd1 vccd1 _12125_/X
+ sky130_fd_sc_hd__o211a_1
X_12056_ hold2564/X hold2722/X _12056_/S vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11007_ _11542_/A _11536_/A _11623_/A _11537_/B vssd1 vssd1 vccd1 vccd1 _11010_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13218__S _13220_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08270__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08478__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ hold819/X hold827/X hold1533/X hold2035/X _12964_/S0 _13068_/A1 vssd1 vssd1
+ vccd1 vccd1 _12958_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08478__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__B1 _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11909_ _13664_/A1 hold1117/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11909_/X sky130_fd_sc_hd__mux2_1
X_12889_ _14289_/Q _14225_/Q hold645/A _14479_/Q _13066_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12889_/X sky130_fd_sc_hd__mux4_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14628_ _15365_/CLK _14628_/D vssd1 vssd1 vccd1 vccd1 _14628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09978__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09978__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ _15429_/CLK hold276/X vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11412__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11785__A1 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _13736_/A1 hold1941/X _07112_/S vssd1 vssd1 vccd1 vccd1 _07100_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08080_ _08080_/A _08080_/B _08080_/C vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__and3_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08650__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07031_ hold663/X _13669_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 hold664/A sky130_fd_sc_hd__mux2_1
XANTENNA__13189__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09386__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10606__A _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__B _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08982_ _08989_/A _08979_/X _08981_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08983_/B
+ sky130_fd_sc_hd__o211a_1
Xhold2704 _14837_/Q vssd1 vssd1 vccd1 vccd1 hold2704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2715 _11102_/Y vssd1 vssd1 vccd1 vccd1 _13402_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _14784_/Q hold939/A hold923/A _14720_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07934_/B sky130_fd_sc_hd__mux4_1
Xhold2726 _15178_/Q vssd1 vssd1 vccd1 vccd1 hold2726/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13636__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2737 _15189_/Q vssd1 vssd1 vccd1 vccd1 hold2737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2748 _15185_/Q vssd1 vssd1 vccd1 vccd1 hold2748/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2759 _15172_/Q vssd1 vssd1 vccd1 vccd1 hold2759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10341__A _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _14084_/Q _14083_/Q _14085_/Q vssd1 vssd1 vccd1 vccd1 _07864_/X sky130_fd_sc_hd__or3_1
XANTENNA__12032__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10512__A2 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _09602_/A _09602_/B _09601_/C _09601_/D vssd1 vssd1 vccd1 vccd1 _09603_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__07126__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10698__D _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07795_ hold1415/X _13700_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 _07795_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11871__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09534_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09534_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_211_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13462__A1 _12288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12896__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10276__A1 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09130__A2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09464_/B _09464_/C _09464_/A vssd1 vssd1 vccd1 vccd1 _09465_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10276__B2 _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout532_A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11172__A _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08416_ _08512_/A _08415_/C _08415_/A vssd1 vssd1 vccd1 vccd1 _08418_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09396_ _10351_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _09398_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_163_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12648__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__A1 _14942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09513__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _08347_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07796__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08278_ _08877_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08278_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07229_ _11606_/A _10304_/D vssd1 vssd1 vccd1 vccd1 _07230_/B sky130_fd_sc_hd__or2_1
XFILLER_0_46_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10516__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ _09514_/A _10239_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _10240_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07827__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _10172_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10171_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13930_ _14754_/CLK _13930_/D vssd1 vssd1 vccd1 vccd1 _13930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07036__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _15458_/CLK hold872/X vssd1 vssd1 vccd1 vccd1 hold871/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11781__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12812_ _06942_/A _12809_/X _12811_/X vssd1 vssd1 vccd1 vccd1 _12812_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_202_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13792_ _06903_/A _13792_/A2 _11693_/X _07475_/B vssd1 vssd1 vccd1 vccd1 _15350_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08656__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_70_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _12749_/S1 _12740_/X _12742_/X vssd1 vssd1 vccd1 vccd1 _12743_/X sky130_fd_sc_hd__a21o_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08880__A1 _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ _13876_/Q _14004_/Q _13844_/Q _13812_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12639__S0 _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14413_ _15446_/CLK hold476/X vssd1 vssd1 vccd1 vccd1 hold475/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _11409_/A _11588_/B _11410_/A _11408_/B vssd1 vssd1 vccd1 vccd1 _11626_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09504__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15393_ _15434_/CLK _15393_/D vssd1 vssd1 vccd1 vccd1 _15393_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12413__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_85_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14344_ _15191_/CLK _14344_/D vssd1 vssd1 vccd1 vccd1 _14344_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08632__A1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ _11620_/A _11586_/B _11376_/A _11374_/B vssd1 vssd1 vccd1 vccd1 _11558_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10507_ _10507_/A _11333_/B _11614_/B _11586_/B vssd1 vssd1 vccd1 vccd1 _10510_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _15045_/CLK _14275_/D vssd1 vssd1 vccd1 vccd1 _14275_/Q sky130_fd_sc_hd__dfxtp_1
X_11487_ _14454_/Q _11486_/B _11486_/Y _07390_/A vssd1 vssd1 vccd1 vccd1 _11487_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10426__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13064__S0 _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13226_ hold1171/X _13738_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10438_ _10351_/A _15221_/Q _10352_/A _10349_/Y vssd1 vssd1 vccd1 vccd1 _10558_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11956__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13389_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _15022_/D sky130_fd_sc_hd__nor2_1
X_10369_ _10191_/X _10193_/Y _10367_/X _10368_/Y vssd1 vssd1 vccd1 vccd1 _10373_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_143_clk_A clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__A2 _10741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ _14994_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12108_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_109_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13456__B _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _06943_/A _13083_/X _13087_/X hold2774/X vssd1 vssd1 vccd1 vccd1 _13095_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_23_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _12059_/A _12039_/B vssd1 vssd1 vccd1 vccd1 _14832_/D sky130_fd_sc_hd__and2_1
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_158_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11407__D _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13472__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07580_ _13719_/A1 hold1637/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07580_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_38_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10258__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13191__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2497_A _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A _14984_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _09250_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08201_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09181_ _09177_/X _09179_/Y _09047_/B _09049_/B vssd1 vssd1 vccd1 vccd1 _09181_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11302__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14581__CLK _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _08564_/A1 _08125_/Y _08127_/Y _08129_/Y _08131_/Y vssd1 vssd1 vccd1 vccd1
+ _08132_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10430__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08063_ _08201_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08063_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07014_ hold755/X _13652_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 hold756/A sky130_fd_sc_hd__mux2_1
XANTENNA__07348__C _15353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12183__A1 hold2555/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12551__A _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2501 _15155_/Q vssd1 vssd1 vccd1 vccd1 hold2501/X sky130_fd_sc_hd__dlygate4sd3_1
X_08965_ _09346_/B _08966_/C _08966_/A vssd1 vssd1 vccd1 vccd1 _08965_/X sky130_fd_sc_hd__o21a_1
Xhold2512 _12069_/X vssd1 vssd1 vccd1 vccd1 _14846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2523 _14876_/Q vssd1 vssd1 vccd1 vccd1 hold2523/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12270__B _12270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_A _07862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2534 hold2848/X vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__buf_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1800 _11944_/X vssd1 vssd1 vccd1 vccd1 _14764_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2545 _13465_/X vssd1 vssd1 vccd1 vccd1 _15226_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07916_ _13342_/A _07915_/B _07908_/X vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__a21o_1
Xhold2556 _12183_/X vssd1 vssd1 vccd1 vccd1 _14902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1811 _14120_/Q vssd1 vssd1 vccd1 vccd1 hold1811/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1822 _07661_/X vssd1 vssd1 vccd1 vccd1 _14282_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08896_ _09136_/A _09866_/B _08895_/C _08895_/D vssd1 vssd1 vccd1 vccd1 _08896_/X
+ sky130_fd_sc_hd__a22o_1
Xhold2567 _15314_/Q vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__clkbuf_2
Xhold2578 _14432_/Q vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__buf_1
Xhold1833 _14408_/Q vssd1 vssd1 vccd1 vccd1 hold1833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2589 _08526_/Y vssd1 vssd1 vccd1 vccd1 hold2589/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1844 _13697_/X vssd1 vssd1 vccd1 vccd1 _15403_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09860__A _09860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1855 _13981_/Q vssd1 vssd1 vccd1 vccd1 hold1855/X sky130_fd_sc_hd__dlygate4sd3_1
X_07847_ hold11/A hold15/A hold17/A hold19/A vssd1 vssd1 vccd1 vccd1 _07847_/X sky130_fd_sc_hd__or4_1
Xhold1866 _07791_/X vssd1 vssd1 vccd1 vccd1 _14406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1877 _14547_/Q vssd1 vssd1 vccd1 vccd1 hold1877/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13382__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1888 _07189_/X vssd1 vssd1 vccd1 vccd1 _13996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1899 _13969_/Q vssd1 vssd1 vccd1 vccd1 hold1899/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10592__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08476__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _13716_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07778_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09517_ _10430_/B1 _09510_/Y _09512_/Y _09514_/Y _09516_/Y vssd1 vssd1 vccd1 vccd1
+ _09517_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11614__B _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _09449_/A _09449_/B _09449_/C vssd1 vssd1 vccd1 vccd1 _09591_/A sky130_fd_sc_hd__o21a_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11333__C _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09379_ _13669_/A1 _11514_/A2 _11514_/B1 _13190_/B _09377_/Y vssd1 vssd1 vccd1 vccd1
+ _09379_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12726__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11410_ _11410_/A _11410_/B vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12390_ hold381/X _14109_/Q _12460_/S vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10421__A1 _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _11341_/A _11341_/B vssd1 vssd1 vccd1 vccd1 _11343_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_132_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08090__A2 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__S0 _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ _15348_/CLK _14060_/D vssd1 vssd1 vccd1 vccd1 _14060_/Q sky130_fd_sc_hd__dfxtp_1
X_11272_ _11273_/A _11273_/B _11273_/C vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_63_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11776__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _13092_/A1 _13010_/X _13100_/S0 vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__a21o_1
X_10223_ _07302_/B _10077_/B _07320_/D vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07555__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _10154_/A _10154_/B _10154_/C vssd1 vssd1 vccd1 vccd1 _10156_/B sky130_fd_sc_hd__and3_2
X_14962_ _14971_/CLK _14962_/D vssd1 vssd1 vccd1 vccd1 _14962_/Q sky130_fd_sc_hd__dfxtp_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ _14446_/Q _13586_/B _10081_/Y hold2502/X _13797_/C1 vssd1 vssd1 vccd1 vccd1
+ _10085_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10488__A1 _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13913_ _15446_/CLK _13913_/D vssd1 vssd1 vccd1 vccd1 _13913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14893_ _14989_/CLK _14893_/D vssd1 vssd1 vccd1 vccd1 _14893_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11227__D _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13844_ _14731_/CLK _13844_/D vssd1 vssd1 vccd1 vccd1 _13844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08386__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11437__B1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13775_ hold217/X vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10987_ _11594_/A _11605_/B _10987_/C _10987_/D vssd1 vssd1 vccd1 vccd1 _10987_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_58_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12726_ _12951_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _12727_/C sky130_fd_sc_hd__or2_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15445_ _15445_/CLK hold428/X vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12657_ _13150_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _14954_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13231__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _11608_/A _11608_/B vssd1 vssd1 vccd1 vccd1 _11609_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10099__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08605__A1 _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15376_ _15376_/CLK _15376_/D vssd1 vssd1 vccd1 vccd1 _15376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12588_ _12642_/B1 _12583_/X _12587_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12595_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09802__B1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12355__B _12379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10412__A1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14327_ _15458_/CLK hold532/X vssd1 vssd1 vccd1 vccd1 hold531/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ _11539_/A _11539_/B vssd1 vssd1 vccd1 vccd1 _11540_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold407 hold407/A vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold418 hold418/A vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09945__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14258_ _15093_/CLK _14258_/D vssd1 vssd1 vccd1 vccd1 _14258_/Q sky130_fd_sc_hd__dfxtp_1
Xhold429 hold429/A vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12165__A1 hold2471/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ hold1097/X _13655_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__mux2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _15188_/CLK hold140/X vssd1 vssd1 vccd1 vccd1 _14189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07465__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13186__B _13186_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2412_A _14068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _08750_/X sky130_fd_sc_hd__or2_1
Xhold1107 _13870_/Q vssd1 vssd1 vccd1 vccd1 hold1107/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _11909_/X vssd1 vssd1 vccd1 vccd1 _14730_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08995__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1129 _14392_/Q vssd1 vssd1 vccd1 vccd1 hold1129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07701_ hold335/X _13674_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold336/A sky130_fd_sc_hd__mux2_1
X_08681_ _08592_/A _08591_/B _08591_/A vssd1 vssd1 vccd1 vccd1 _08694_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__08767__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07632_ hold1081/X _13738_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07632_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_178_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2781_A _15193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _13396_/A hold191/X vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__and2_1
X_09302_ _10185_/A _09709_/B _09301_/C _09400_/A vssd1 vssd1 vccd1 vccd1 _09303_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11153__C _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__A1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ hold1083/X _13700_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07494_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09233_ _14347_/Q _14251_/Q hold977/A _14123_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09234_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12928__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08743__B _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09164_ _09164_/A _09979_/D _09165_/A vssd1 vssd1 vccd1 vccd1 _09164_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12265__B _13416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08115_ hold187/A hold333/A _14595_/Q _13964_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08115_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_161_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09095_ hold283/A _14314_/Q hold585/A _13974_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09095_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08072__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08046_ _13554_/B _08046_/B _08046_/C vssd1 vssd1 vccd1 vccd1 _08046_/X sky130_fd_sc_hd__or3_1
XFILLER_0_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold930 hold930/A vssd1 vssd1 vccd1 vccd1 hold930/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold941 hold941/A vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 hold952/A vssd1 vssd1 vccd1 vccd1 hold952/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13377__A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 hold963/A vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12281__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 hold974/A vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 hold996/A vssd1 vssd1 vccd1 vccd1 hold996/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ _09997_/A _09997_/B _09997_/C vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__nand3_2
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout864_A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2320 _12133_/X vssd1 vssd1 vccd1 vccd1 _14877_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2331 _15342_/Q vssd1 vssd1 vccd1 vccd1 hold2331/X sky130_fd_sc_hd__buf_1
XFILLER_0_157_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _08948_/A _08948_/B _08948_/C vssd1 vssd1 vccd1 vccd1 _08997_/A sky130_fd_sc_hd__nand3_2
Xhold2342 hold2840/X vssd1 vssd1 vccd1 vccd1 _07432_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2353 _12169_/X vssd1 vssd1 vccd1 vccd1 _14895_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2364 _14028_/Q vssd1 vssd1 vccd1 vccd1 _06923_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1630 _11957_/X vssd1 vssd1 vccd1 vccd1 _14777_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2375 _15035_/Q vssd1 vssd1 vccd1 vccd1 _07575_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1641 _14556_/Q vssd1 vssd1 vccd1 vccd1 hold1641/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2386 _14062_/Q vssd1 vssd1 vccd1 vccd1 _06921_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1652 _11708_/X vssd1 vssd1 vccd1 vccd1 _14504_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08879_ _08873_/A _08878_/X _08880_/A1 vssd1 vssd1 vccd1 vccd1 _08879_/Y sky130_fd_sc_hd__o21ai_1
Xhold2397 _13565_/X vssd1 vssd1 vccd1 vccd1 _15308_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1663 _13980_/Q vssd1 vssd1 vccd1 vccd1 hold1663/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08918__B _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1674 _11856_/X vssd1 vssd1 vccd1 vccd1 _14679_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _11098_/B _10909_/X _10726_/Y _10730_/A vssd1 vssd1 vccd1 vccd1 _10910_/X
+ sky130_fd_sc_hd__o211a_1
Xhold1685 _14636_/Q vssd1 vssd1 vccd1 vccd1 hold1685/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12220__S _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1696 _07583_/X vssd1 vssd1 vccd1 vccd1 _14207_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13408__A1 _12261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ hold1037/X _13711_/A1 _11893_/S vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _11409_/A _11390_/A _10840_/C _10840_/D vssd1 vssd1 vccd1 vccd1 _10841_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_168_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07099__A0 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _14436_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10772_ _15417_/Q hold869/A _14712_/Q hold773/A _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10772_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_137_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12631__A2 _13152_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _12692_/A1 _12510_/X _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12511_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ _13491_/A hold53/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__and2_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ _15258_/CLK _15230_/D vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _12642_/A1 _12441_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12442_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15189__D _15189_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _15296_/CLK _15161_/D vssd1 vssd1 vccd1 vccd1 _15161_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07269__B _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12890__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12373_ hold763/A _14719_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12373_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14112_ _15428_/CLK _14112_/D vssd1 vssd1 vccd1 vccd1 _14112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _07240_/B _11323_/X _07328_/A vssd1 vssd1 vccd1 vccd1 _11324_/X sky130_fd_sc_hd__a21o_1
X_15092_ _15408_/CLK _15092_/D vssd1 vssd1 vccd1 vccd1 _15092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12147__A1 hold2634/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13287__A _13287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14043_ _15293_/CLK hold106/X vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
X_11255_ _11254_/B _11254_/C _11254_/A vssd1 vssd1 vccd1 vccd1 _11255_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08446__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12242__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _10206_/A _10206_/B _10206_/C _10206_/D vssd1 vssd1 vccd1 vccd1 _10206_/X
+ sky130_fd_sc_hd__or4_4
XANTENNA__07285__A _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10253__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _11220_/A vssd1 vssd1 vccd1 vccd1 _11455_/A sky130_fd_sc_hd__inv_2
XFILLER_0_24_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _10024_/C _10023_/Y _10135_/Y _10136_/X vssd1 vssd1 vccd1 vccd1 _10137_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13647__A1 _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10142__C _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09946__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ _10064_/X _10066_/Y _09903_/Y _09905_/X vssd1 vssd1 vccd1 vccd1 _10263_/B
+ sky130_fd_sc_hd__o211a_1
X_14945_ _15214_/CLK _14945_/D vssd1 vssd1 vccd1 vccd1 _14945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13226__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ _14876_/CLK _14876_/D vssd1 vssd1 vccd1 vccd1 _14876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13827_ _15458_/CLK _13827_/D vssd1 vssd1 vccd1 vccd1 _13827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13750__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13758_ hold275/X vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ hold395/X _13910_/Q _12791_/S vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09659__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13689_ hold1529/X _13689_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12366__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15428_ _15428_/CLK _15428_/D vssd1 vssd1 vccd1 vccd1 _15428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12386__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15359_ _15428_/CLK hold884/X vssd1 vssd1 vccd1 vccd1 hold883/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13197__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _09778_/A _09930_/A _09774_/A vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 _13690_/A1 vssd1 vssd1 vccd1 vccd1 _13657_/A1 sky130_fd_sc_hd__clkbuf_4
X_09851_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__nand2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__A0 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 _15038_/Q vssd1 vssd1 vccd1 vccd1 _13652_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__11429__B _14970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 _10283_/C vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__08988__S1 _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _14954_/Q vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__buf_4
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__xnor2_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _15153_/Q _09925_/A2 _13590_/B vssd1 vssd1 vccd1 vccd1 _09782_/Y sky130_fd_sc_hd__a21oi_1
X_06994_ _13666_/A1 hold1551/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06994_/X sky130_fd_sc_hd__mux2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08571_/A _08571_/B _08628_/A _08734_/A _08629_/A vssd1 vssd1 vccd1 vccd1
+ _08841_/B sky130_fd_sc_hd__o311ai_4
XANTENNA__07923__A _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08981_/A _08663_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08664_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07134__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07615_ hold1517/X _13721_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07615_/X sky130_fd_sc_hd__mux2_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _09164_/A _09858_/C vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout445_A _07389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07546_ _13386_/A hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__and2_1
XFILLER_0_152_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10624__A1 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout612_A _15207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__A2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ _11928_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07477_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12276__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _09217_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12377__A1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ _09146_/B _09146_/C _09146_/A vssd1 vssd1 vccd1 vccd1 _09148_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09242__B2 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10927__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ _11640_/B1 _09074_/X _09075_/X _09077_/Y vssd1 vssd1 vccd1 vccd1 _13389_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _07283_/A _07951_/B _07283_/B vssd1 vssd1 vccd1 vccd1 _08029_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_60_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold760 hold760/A vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 hold771/A vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 hold782/A vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _11526_/A _11333_/B _15221_/Q _15222_/Q vssd1 vssd1 vccd1 vccd1 _11229_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08979__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 hold793/A vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2150 _13513_/X vssd1 vssd1 vccd1 vccd1 _15271_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2161 _15261_/Q vssd1 vssd1 vccd1 vccd1 hold2161/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2172 _11676_/X vssd1 vssd1 vccd1 vccd1 _14479_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2183 _13942_/Q vssd1 vssd1 vccd1 vccd1 hold2183/X sky130_fd_sc_hd__dlygate4sd3_1
X_12991_ hold735/X hold903/X _12991_/S vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__mux2_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2194 _07005_/X vssd1 vssd1 vccd1 vccd1 _13824_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1460 _07157_/X vssd1 vssd1 vccd1 vccd1 _13965_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14730_ _15369_/CLK _14730_/D vssd1 vssd1 vccd1 vccd1 _14730_/Q sky130_fd_sc_hd__dfxtp_1
X_11942_ _13730_/A1 hold2215/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11942_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1471 _14789_/Q vssd1 vssd1 vccd1 vccd1 hold1471/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1482 _07003_/X vssd1 vssd1 vccd1 vccd1 _13822_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 _14626_/Q vssd1 vssd1 vccd1 vccd1 hold1493/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07044__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14661_ _15435_/CLK _14661_/D vssd1 vssd1 vccd1 vccd1 _14661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12885__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ hold429/X _13727_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold430/A sky130_fd_sc_hd__mux2_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13612_ _07429_/A _13625_/C _13611_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15333_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10824_ _11620_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _10825_/B sky130_fd_sc_hd__nand2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08808__A1 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _15072_/CLK hold972/X vssd1 vssd1 vccd1 vccd1 hold971/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12604__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13543_ _07974_/A _13591_/A2 _13542_/X _13541_/A vssd1 vssd1 vccd1 vccd1 _13543_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ _11104_/A _12286_/B _10750_/Y _10754_/X vssd1 vssd1 vccd1 vccd1 _10755_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13474_ _13481_/A _13474_/B vssd1 vssd1 vccd1 vccd1 _15233_/D sky130_fd_sc_hd__and2_2
XFILLER_0_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10686_ _10686_/A _10686_/B vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__or2_1
XFILLER_0_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _15427_/CLK _15213_/D vssd1 vssd1 vccd1 vccd1 _15213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ _12421_/X _12422_/X _12424_/X _12423_/X _12644_/A1 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12426_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15144_ _15305_/CLK _15144_/D vssd1 vssd1 vccd1 vccd1 _15144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09784__A2 _13446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _13173_/B _12953_/B1 _12354_/X _13718_/A1 _12355_/X vssd1 vssd1 vccd1 vccd1
+ _12356_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput309 _14870_/Q vssd1 vssd1 vccd1 vccd1 out1[25] sky130_fd_sc_hd__buf_12
XANTENNA__06912__A _15341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11507_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15075_ _15299_/CLK _15075_/D vssd1 vssd1 vccd1 vccd1 _15075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12287_ _13171_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _14936_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12215__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14026_ _15348_/CLK hold272/X vssd1 vssd1 vccd1 vccd1 _14026_/Q sky130_fd_sc_hd__dfxtp_1
X_11238_ _11567_/A _15226_/Q _11239_/A vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__and3_1
XANTENNA__11964__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _11169_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11177_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_207_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__B _13464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14928_ _15251_/CLK _14928_/D vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14859_ _15004_/CLK _14859_/D vssd1 vssd1 vccd1 vccd1 _14859_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12056__A0 hold2564/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07400_ hold573/X _07448_/B vssd1 vssd1 vccd1 vccd1 hold574/A sky130_fd_sc_hd__and2_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _08380_/A _08380_/B vssd1 vssd1 vccd1 vccd1 _08429_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08574__A _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07331_ _07221_/A _07323_/A _07321_/Y _07330_/X vssd1 vssd1 vccd1 vccd1 _12221_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12096__A _14988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07262_ _15227_/Q _14971_/Q vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ _09001_/A _09127_/A vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_155_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold2744_A _15179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07193_ hold1825/X _13661_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 _07193_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11319__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07129__S _07131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ _09903_/A vssd1 vssd1 vccd1 vccd1 _09903_/Y sky130_fd_sc_hd__inv_2
Xfanout503 _06942_/Y vssd1 vssd1 vccd1 vccd1 _12692_/A1 sky130_fd_sc_hd__buf_6
Xfanout514 _10252_/A vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__buf_6
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout525 _10255_/A1 vssd1 vssd1 vccd1 vccd1 _10430_/B1 sky130_fd_sc_hd__buf_6
XANTENNA__07538__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 _11507_/A vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__11874__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _07677_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ _09833_/B _09833_/C _09833_/A vssd1 vssd1 vccd1 vccd1 _09834_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12531__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _10087_/S1 vssd1 vssd1 vccd1 vccd1 _09239_/S1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10768__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 _08763_/S0 vssd1 vssd1 vccd1 vccd1 _08130_/S0 sky130_fd_sc_hd__buf_8
Xfanout569 _10425_/S0 vssd1 vssd1 vccd1 vccd1 _10429_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_193_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09765_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__and2_1
XANTENNA__13374__B _13374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06977_ _07875_/B _07114_/B vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__or2_2
XANTENNA__12819__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_A _08275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ _08717_/A _08717_/B _08717_/C vssd1 vssd1 vccd1 vccd1 _08716_/X sky130_fd_sc_hd__and3_1
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09696_ _09745_/A vssd1 vssd1 vccd1 vccd1 _09696_/Y sky130_fd_sc_hd__inv_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _08750_/A _08856_/C vssd1 vssd1 vccd1 vccd1 _08647_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout827_A _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10940__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07799__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13390__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08901_/A _09866_/B _08577_/C vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__a21oi_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ hold1115/X _13700_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 _07529_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10540_ _10537_/X _10538_/Y _10364_/X _10366_/Y vssd1 vssd1 vccd1 vccd1 _10541_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10471_ _11620_/A _11378_/C vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_161_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11060__D _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13753__A2_N _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _12243_/A _12210_/B vssd1 vssd1 vccd1 vccd1 _12210_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07828__A _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ _13397_/A _13190_/B vssd1 vssd1 vccd1 vccd1 _15055_/D sky130_fd_sc_hd__and2_1
XFILLER_0_121_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ hold2628/X _12173_/A2 _12140_/X _13486_/A vssd1 vssd1 vccd1 vccd1 _12141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07039__S _07044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ _14976_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12072_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold590 hold590/A vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11784__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _11022_/B _11022_/C _11022_/A vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_60_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07563__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13078__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__B _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _13888_/Q _14016_/Q _13856_/Q _13824_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12974_/X sky130_fd_sc_hd__mux4_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1290 _11869_/X vssd1 vssd1 vccd1 vccd1 _14691_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _15455_/CLK hold732/X vssd1 vssd1 vccd1 vccd1 hold731/A sky130_fd_sc_hd__dfxtp_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _13680_/A1 hold1087/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__mux2_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__A0 hold2593/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13504__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _15408_/CLK hold848/X vssd1 vssd1 vccd1 vccd1 hold847/A sky130_fd_sc_hd__dfxtp_1
X_11856_ hold1673/X _13743_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__mux2_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _11573_/A _11605_/B _10807_/C _10807_/D vssd1 vssd1 vccd1 vccd1 _10807_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_0_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14575_ _15410_/CLK hold240/X vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11787_ hold1123/X _13674_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 _11787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09002__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10738_ _10958_/A _10737_/X _11473_/A vssd1 vssd1 vccd1 vccd1 _10738_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13526_ _13740_/A1 hold1731/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13526_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11959__S _11959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ _10568_/B _13466_/A _13456_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 _15222_/D
+ sky130_fd_sc_hd__o211a_1
X_10669_ _10669_/A vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ hold1643/X _14529_/Q hold671/X hold1881/X _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12408_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_140_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13388_ _13393_/A _13388_/B vssd1 vssd1 vccd1 vccd1 _15179_/D sky130_fd_sc_hd__and2_1
XFILLER_0_140_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12761__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15127_ _15127_/CLK _15127_/D vssd1 vssd1 vccd1 vccd1 _15127_/Q sky130_fd_sc_hd__dfxtp_1
X_12339_ _12335_/X _12336_/X _12338_/X _12337_/X _12366_/A _06944_/A vssd1 vssd1 vccd1
+ vccd1 _12339_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15058_ _15443_/CLK _15058_/D vssd1 vssd1 vccd1 vccd1 _15058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12513__A1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ _15444_/CLK _14009_/D vssd1 vssd1 vccd1 vccd1 _14009_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10314__D _14957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13475__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _07879_/A _12379_/B _07900_/A vssd1 vssd1 vccd1 vccd1 _07899_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__13194__B _13194_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09550_ _09549_/B _09549_/C _09549_/A vssd1 vssd1 vccd1 vccd1 _09550_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_211_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08501_ _08500_/B _08500_/C _08500_/A vssd1 vssd1 vccd1 vccd1 _08502_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09481_ _09481_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09481_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_hold2694_A _15167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _07900_/B _13383_/B _08376_/X vssd1 vssd1 vccd1 vccd1 _13424_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2861_A _15345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08363_ _12241_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08363_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12675__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07314_ _09437_/A _11351_/B vssd1 vssd1 vccd1 vccd1 _08338_/C sky130_fd_sc_hd__or2_1
X_08294_ _08776_/A _08926_/A _08294_/C _08294_/D vssd1 vssd1 vccd1 vccd1 _08401_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11869__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ _09864_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _08528_/D sky130_fd_sc_hd__or2_1
XFILLER_0_117_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout408_A _07149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07176_ hold2765/A hold1779/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07176_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12273__B _12273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09863__A _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13385__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__A1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09074__S _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 _07903_/Y vssd1 vssd1 vccd1 vccd1 _13750_/A sky130_fd_sc_hd__clkbuf_8
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__xor2_1
Xfanout377 _12325_/B vssd1 vssd1 vccd1 vccd1 _13104_/A2 sky130_fd_sc_hd__buf_6
Xfanout388 _11696_/Y vssd1 vssd1 vccd1 vccd1 _11728_/S sky130_fd_sc_hd__buf_12
XFILLER_0_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10521__B _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _07577_/Y vssd1 vssd1 vccd1 vccd1 _07593_/S sky130_fd_sc_hd__buf_12
XFILLER_0_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07931__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09359__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _09744_/Y _09746_/X _09601_/C _09602_/X vssd1 vssd1 vccd1 vccd1 _09748_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13465__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12363__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A _09679_/B _09824_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__nand3_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__B _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ hold725/X _13664_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold726/A sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12690_ hold747/X hold857/A _12741_/S vssd1 vssd1 vccd1 vccd1 _12690_/X sky130_fd_sc_hd__mux2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11641_ _11515_/Y _11516_/X _11639_/X _11640_/X vssd1 vssd1 vccd1 vccd1 _11641_/X
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__11352__B _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11243__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14360_ _15068_/CLK hold658/X vssd1 vssd1 vccd1 vccd1 hold657/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11243__B2 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _11572_/A _11572_/B vssd1 vssd1 vccd1 vccd1 _11583_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08644__C1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13311_ _13317_/A _13311_/B vssd1 vssd1 vccd1 vccd1 _15123_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11779__S _11779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10523_ _10311_/A _10310_/B _10308_/X vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__a21o_1
Xinput19 dmemresp_rdata[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
X_14291_ _15415_/CLK _14291_/D vssd1 vssd1 vccd1 vccd1 _14291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ fanout6/X fanout4/X vssd1 vssd1 vccd1 vccd1 fanout2/A sky130_fd_sc_hd__nor2_1
XFILLER_0_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07558__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _10455_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _10454_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12743__A1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13173_ _13481_/A _13173_/B vssd1 vssd1 vccd1 vccd1 _15038_/D sky130_fd_sc_hd__and2_1
X_10385_ _10382_/Y _10383_/X _10201_/X _10204_/Y vssd1 vssd1 vccd1 vccd1 _10387_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10754__B1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _15002_/Q _12126_/B _12126_/C _12124_/D vssd1 vssd1 vccd1 vccd1 _12124_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__09773__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ _12059_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _14840_/D sky130_fd_sc_hd__and2_1
X_11006_ _11542_/A _11536_/A _11623_/A _11537_/B vssd1 vssd1 vccd1 vccd1 _11006_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__08270__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__B1 _13375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08478__A2 _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _13171_/A _12957_/B vssd1 vssd1 vccd1 vccd1 _14966_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09675__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13234__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ _13663_/A1 hold2087/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11908_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12888_ _12917_/B1 _12883_/X _12887_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12895_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _15299_/CLK hold996/X vssd1 vssd1 vccd1 vccd1 hold995/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11839_ hold1303/X _15046_/Q _11845_/S vssd1 vssd1 vccd1 vccd1 _11839_/X sky130_fd_sc_hd__mux2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09978__A2 _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12431__B1 _13144_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ _15364_/CLK hold252/X vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13657_/A1 hold1885/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ _15348_/CLK _14489_/D vssd1 vssd1 vccd1 vccd1 _14489_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07030_ hold1999/X _13668_/A1 _07044_/S vssd1 vssd1 vccd1 vccd1 _07030_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09386__C _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10606__B _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2442_A _11474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08981_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _08981_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2705 _14835_/Q vssd1 vssd1 vccd1 vccd1 hold2705/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold2707_A _10741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ _15361_/Q _15264_/Q hold935/A _14365_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _07932_/X sky130_fd_sc_hd__mux4_1
Xhold2716 _14839_/Q vssd1 vssd1 vccd1 vccd1 hold2716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2727 _15187_/Q vssd1 vssd1 vccd1 vccd1 hold2727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2738 _15182_/Q vssd1 vssd1 vccd1 vccd1 hold2738/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07955__A1_N _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2749 _15061_/Q vssd1 vssd1 vccd1 vccd1 hold2749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07863_ _14084_/Q _14083_/Q _14085_/Q vssd1 vssd1 vccd1 vccd1 _07863_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_208_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10341__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11170__B1 _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09602_ _09602_/A _09602_/B _09601_/C _09601_/D vssd1 vssd1 vccd1 vccd1 _09602_/X
+ sky130_fd_sc_hd__or4bb_2
X_07794_ hold747/X _13732_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold748/A sky130_fd_sc_hd__mux2_1
X_09533_ _09533_/A _09533_/B vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12896__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A _12330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _09464_/A _09464_/B _09464_/C vssd1 vssd1 vccd1 vccd1 _09464_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_149_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10276__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12268__B _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07142__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ _08415_/A _08512_/A _08415_/C vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11172__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09395_ _09395_/A _09395_/B vssd1 vssd1 vccd1 vccd1 _09398_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout525_A _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12648__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ _08344_/Y _08346_/B vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09969__A2 _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08277_ hold379/A hold495/A _14146_/Q _14464_/Q _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08278_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12284__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10984__B1 _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07228_ _11606_/A _10304_/D vssd1 vssd1 vccd1 vccd1 _07230_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout894_A input161/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10516__B _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ _13512_/A0 hold1901/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07827__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ _10170_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__or2_2
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08002__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13860_ _15384_/CLK _13860_/D vssd1 vssd1 vccd1 vccd1 _13860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12336__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ _12917_/A1 _12810_/X _12844_/A1 vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13562__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13791_ _06904_/A _13792_/A2 _11691_/X _07475_/B vssd1 vssd1 vccd1 vccd1 _15349_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13453__A2 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12917_/A1 _12741_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12742_/X sky130_fd_sc_hd__a21o_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__B1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07052__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ hold231/A _14312_/Q _14603_/Q _13972_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12673_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_210_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__S1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11624_ _11622_/X _11392_/B _11624_/S vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__mux2_1
X_14412_ _15410_/CLK hold584/X vssd1 vssd1 vccd1 vccd1 hold583/A sky130_fd_sc_hd__dfxtp_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15392_ _15392_/CLK _15392_/D vssd1 vssd1 vccd1 vccd1 _15392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ _11555_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14343_ _15405_/CLK hold990/X vssd1 vssd1 vccd1 vccd1 hold989/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07288__A _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ _10502_/Y _10503_/X _10295_/Y _10332_/X vssd1 vssd1 vccd1 vccd1 _10548_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_107_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14274_ _14954_/CLK hold380/X vssd1 vssd1 vccd1 vccd1 hold379/A sky130_fd_sc_hd__dfxtp_1
X_11486_ _14454_/Q _11486_/B vssd1 vssd1 vccd1 vccd1 _11486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ hold307/X _13671_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__mux2_1
X_10437_ _10600_/A _07280_/B _10262_/X _11640_/B1 vssd1 vssd1 vccd1 vccd1 _10437_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08396__A1 _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _13389_/A _13156_/B vssd1 vssd1 vccd1 vccd1 _15021_/D sky130_fd_sc_hd__nor2_1
X_10368_ _10364_/X _10365_/Y _10189_/B _10191_/B vssd1 vssd1 vccd1 vccd1 _10368_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ hold2475/X _12129_/A2 _12106_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12107_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13229__S _13236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13099_/S1 _13084_/X _13086_/X vssd1 vssd1 vccd1 vccd1 _13087_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_209_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10299_ _10827_/D _10297_/X _10298_/X vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09008__A _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ hold2593/X hold2712/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12039_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12575__S0 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__B1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13989_ _15292_/CLK _13989_/D vssd1 vssd1 vccd1 vccd1 _13989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_181_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08200_ _14660_/Q _13933_/Q _15434_/Q _13901_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08201_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_34_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ _09047_/B _09049_/B _09177_/X _09179_/Y vssd1 vssd1 vccd1 vccd1 _09180_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__09678__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08582__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12955__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08131_ _08197_/A _08130_/X _08564_/A1 vssd1 vssd1 vccd1 vccd1 _08131_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11302__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__B _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10617__A _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10966__B1 _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08062_ hold503/A _14207_/Q _14143_/Q _14461_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08063_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_114_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07013_ hold1969/X _13651_/A1 _07028_/S vssd1 vssd1 vccd1 vccd1 _07013_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07348__D _15352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2502 _10084_/X vssd1 vssd1 vccd1 vccd1 hold2502/X sky130_fd_sc_hd__dlygate4sd3_1
X_08964_ _08964_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _08966_/C sky130_fd_sc_hd__and2_1
Xhold2513 _14848_/Q vssd1 vssd1 vccd1 vccd1 hold2513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2524 _12129_/X vssd1 vssd1 vccd1 vccd1 _14876_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07137__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2535 _14999_/Q vssd1 vssd1 vccd1 vccd1 hold2535/X sky130_fd_sc_hd__buf_2
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07915_ _07908_/X _07915_/B vssd1 vssd1 vccd1 vccd1 _13342_/B sky130_fd_sc_hd__nand2b_1
Xhold1801 _13816_/Q vssd1 vssd1 vccd1 vccd1 hold1801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2546 _14451_/Q vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08895_ _09136_/A _09866_/B _08895_/C _08895_/D vssd1 vssd1 vccd1 vccd1 _08895_/Y
+ sky130_fd_sc_hd__nand4_1
Xhold2557 _15352_/Q vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__buf_2
Xhold1812 _07492_/X vssd1 vssd1 vccd1 vccd1 _14120_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _13873_/Q vssd1 vssd1 vccd1 vccd1 hold1823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2568 _13577_/X vssd1 vssd1 vccd1 vccd1 _15314_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout475_A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2579 _08351_/X vssd1 vssd1 vccd1 vccd1 _14432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1834 _07793_/X vssd1 vssd1 vccd1 vccd1 _14408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1845 _15273_/Q vssd1 vssd1 vccd1 vccd1 hold1845/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09860__B _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _07846_/A _12308_/B _07846_/C vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10167__A1_N _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1856 _07173_/X vssd1 vssd1 vccd1 vccd1 _13981_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1867 _15376_/Q vssd1 vssd1 vccd1 vccd1 hold1867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1878 _11753_/X vssd1 vssd1 vccd1 vccd1 _14547_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1889 _13869_/Q vssd1 vssd1 vccd1 vccd1 hold1889/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12318__S0 _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13382__B _13382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14909__D _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _13748_/A1 hold1279/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07777_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout642_A _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__A _13168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08476__B _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09516_ _09941_/A _09515_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09516_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09579_/B _09447_/B vssd1 vssd1 vccd1 vccd1 _09449_/C sky130_fd_sc_hd__and2_1
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11333__D _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_172_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _14602_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09378_ hold2703/X input10/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13190_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07600__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ _08329_/A _08329_/B _08329_/C vssd1 vssd1 vccd1 vccd1 _08331_/B sky130_fd_sc_hd__and3_1
XFILLER_0_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10957__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ _11340_/A _15226_/Q vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13046__S1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11271_ _11465_/B _11271_/B vssd1 vssd1 vccd1 vccd1 _11273_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ hold651/X hold1957/X _13041_/S vssd1 vssd1 vccd1 vccd1 _13010_/X sky130_fd_sc_hd__mux2_1
X_10222_ hold2731/X _11283_/S _11640_/B1 vssd1 vssd1 vccd1 vccd1 _10222_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10152_/A _10152_/B _10152_/C vssd1 vssd1 vccd1 vccd1 _10154_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07047__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14961_ _14971_/CLK _14961_/D vssd1 vssd1 vccd1 vccd1 _14961_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10084_ hold2501/X _07812_/A _13590_/B _09934_/Y _10083_/Y vssd1 vssd1 vccd1 vccd1
+ _10084_/X sky130_fd_sc_hd__a2111o_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11792__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ _15445_/CLK _13912_/D vssd1 vssd1 vccd1 vccd1 _13912_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10488__A2 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08667__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ _14989_/CLK _14892_/D vssd1 vssd1 vccd1 vccd1 _14892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08550__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13843_ _15369_/CLK _13843_/D vssd1 vssd1 vccd1 vccd1 _13843_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08386__B _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11437__A1 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11437__B2 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ _11594_/A _11605_/B _10987_/C _10987_/D vssd1 vssd1 vccd1 vccd1 _10986_/X
+ sky130_fd_sc_hd__a22o_1
X_13774_ hold239/X vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__08302__A1 _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12725_ _12721_/X _12722_/X _12724_/X _12723_/X _12844_/A1 _12944_/C1 vssd1 vssd1
+ vccd1 vccd1 _12726_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_163_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_183_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13512__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15444_ _15444_/CLK hold724/X vssd1 vssd1 vccd1 vccd1 hold723/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ _13106_/A1 _13153_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12937__A1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _11607_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__nand2_1
X_15375_ _15375_/CLK hold374/X vssd1 vssd1 vccd1 vccd1 hold373/A sky130_fd_sc_hd__dfxtp_1
X_12587_ _12699_/S1 _12584_/X _12586_/X vssd1 vssd1 vccd1 vccd1 _12587_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10099__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08605__A2 _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09802__A1 _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12355__C _13375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10412__A2 _12284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14326_ _14483_/CLK hold318/X vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__dfxtp_1
X_11538_ _11538_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold408 hold408/A vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11967__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold419 hold419/A vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _11470_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _11469_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14257_ _15196_/CLK _14257_/D vssd1 vssd1 vccd1 vccd1 _14257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12652__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__B1 _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ hold935/X _13654_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 hold936/A sky130_fd_sc_hd__mux2_1
XANTENNA__12796__S0 _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10176__A1 _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188_ _15188_/CLK hold192/X vssd1 vssd1 vccd1 vccd1 _14188_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _13501_/A hold707/X vssd1 vssd1 vccd1 vccd1 hold708/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12548__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _07054_/X vssd1 vssd1 vccd1 vccd1 _13870_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1119 _15448_/Q vssd1 vssd1 vccd1 vccd1 hold1119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07700_ hold559/X _13673_/A1 _07709_/S vssd1 vssd1 vccd1 vccd1 hold560/A sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13483__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ _08816_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _08680_/X sky130_fd_sc_hd__or2_1
XFILLER_0_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08577__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07631_ hold533/X _13737_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 hold534/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13417__A2 _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07562_ _13396_/A hold119/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__and2_1
XFILLER_0_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09301_ _10185_/A _09709_/B _09301_/C _09400_/A vssd1 vssd1 vccd1 vccd1 _09400_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2774_A _14491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07493_ hold857/X _13732_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 hold858/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_154_clk clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _15436_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11153__D _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12827__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09232_ _10246_/A _09232_/B vssd1 vssd1 vccd1 vccd1 _09232_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_173_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12928__A1 _13708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08743__C _08743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09163_ _09164_/A _09979_/D vssd1 vssd1 vccd1 vccd1 _09165_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12928__B2 _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08114_ _14430_/Q _08257_/C vssd1 vssd1 vccd1 vccd1 _08114_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ _09350_/B _09350_/C vssd1 vssd1 vccd1 vccd1 _09094_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11877__S _11877_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ _09494_/A1 _08043_/Y _08044_/X _09925_/A2 hold2583/X vssd1 vssd1 vccd1 vccd1
+ _08045_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_141_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold920 hold920/A vssd1 vssd1 vccd1 vccd1 hold920/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold931 hold931/A vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold942 hold942/A vssd1 vssd1 vccd1 vccd1 hold942/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13377__B _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold953 hold953/A vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 hold964/A vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__B _13448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 hold975/A vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 hold986/A vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 hold997/A vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ _09995_/B _09995_/C _09995_/A vssd1 vssd1 vccd1 vccd1 _09997_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2310 hold2824/X vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__buf_1
XANTENNA__13105__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2321 hold2850/X vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12539__S0 _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2332 _13794_/X vssd1 vssd1 vccd1 vccd1 _15423_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _08944_/Y _08945_/X _08829_/B _08829_/Y vssd1 vssd1 vccd1 vccd1 _08948_/C
+ sky130_fd_sc_hd__a211o_1
Xhold2343 hold2844/X vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__buf_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout857_A _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2354 hold2838/X vssd1 vssd1 vccd1 vccd1 hold2354/X sky130_fd_sc_hd__buf_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2365 _15133_/Q vssd1 vssd1 vccd1 vccd1 hold2365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1620 _07729_/X vssd1 vssd1 vccd1 vccd1 _14348_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13393__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2376 _15040_/Q vssd1 vssd1 vccd1 vccd1 hold2376/X sky130_fd_sc_hd__buf_1
Xhold1631 _14460_/Q vssd1 vssd1 vccd1 vccd1 hold1631/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_84_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2387 hold2836/X vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__buf_1
Xhold1642 _11762_/X vssd1 vssd1 vccd1 vccd1 _14556_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2398 _14860_/Q vssd1 vssd1 vccd1 vccd1 hold2398/X sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ hold909/A hold653/A _14699_/Q _14763_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08878_/X sky130_fd_sc_hd__mux4_1
Xhold1653 _13863_/Q vssd1 vssd1 vccd1 vccd1 hold1653/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1664 _07172_/X vssd1 vssd1 vccd1 vccd1 _13980_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07391__A _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1675 _14347_/Q vssd1 vssd1 vccd1 vccd1 hold1675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ _14268_/Q _14204_/Q _14140_/Q _14458_/Q _12237_/S _12211_/S1 vssd1 vssd1
+ vccd1 vccd1 _07830_/B sky130_fd_sc_hd__mux4_1
Xhold1686 _11812_/X vssd1 vssd1 vccd1 vccd1 _14636_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1697 _14632_/Q vssd1 vssd1 vccd1 vccd1 hold1697/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ _11409_/A _11390_/A _10840_/C _10840_/D vssd1 vssd1 vccd1 vccd1 _11015_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_196_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_99_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _11504_/A _10771_/B vssd1 vssd1 vccd1 vccd1 _10771_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_145_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15453_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_142_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _14661_/Q _13934_/Q _12560_/S vssd1 vssd1 vccd1 vccd1 _12510_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13490_ _13490_/A hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__and2_1
XFILLER_0_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12919__A1 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ hold415/A _14239_/Q _12441_/S vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_22_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10257__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12372_ _14783_/Q _14495_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__mux2_1
X_15160_ _15325_/CLK _15160_/D vssd1 vssd1 vccd1 vccd1 _15160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_157_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ _11285_/A _11285_/B _07240_/A vssd1 vssd1 vccd1 vccd1 _11323_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__11787__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14111_ _15391_/CLK _14111_/D vssd1 vssd1 vccd1 vccd1 _14111_/Q sky130_fd_sc_hd__dfxtp_1
X_15091_ _15441_/CLK hold838/X vssd1 vssd1 vccd1 vccd1 hold837/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07566__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _11254_/A _11254_/B _11254_/C vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__nand3_2
X_14042_ _14042_/CLK _14042_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_37_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08446__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _10201_/X _10202_/Y _09993_/B _09995_/B vssd1 vssd1 vccd1 vccd1 _10206_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__07285__B _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11185_ _10996_/A _10996_/Y _11183_/Y _11184_/X vssd1 vssd1 vccd1 vccd1 _11220_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10253__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10136_ _10306_/A _11168_/A _10135_/C _10135_/D vssd1 vssd1 vccd1 vccd1 _10136_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09781__A _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13647__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13507__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__D _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10067_ _09903_/Y _09905_/X _10064_/X _10066_/Y vssd1 vssd1 vccd1 vccd1 _10266_/B
+ sky130_fd_sc_hd__a211oi_2
X_14944_ _15293_/CLK _14944_/D vssd1 vssd1 vccd1 vccd1 _14944_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09946__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12950__S0 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ _14876_/CLK _14875_/D vssd1 vssd1 vccd1 vccd1 _14875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5__f_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13826_ _15196_/CLK _13826_/D vssd1 vssd1 vccd1 vccd1 _13826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08287__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ hold251/X vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_136_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_168_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _11598_/A _11594_/B _10969_/C _11150_/A vssd1 vssd1 vccd1 vccd1 _11150_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ hold405/X _14541_/Q hold987/A _14765_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12708_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09659__C _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13688_ hold1643/X _13721_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 _13688_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ _15427_/CLK _15427_/D vssd1 vssd1 vccd1 vccd1 _15427_/Q sky130_fd_sc_hd__dfxtp_1
X_12639_ _14279_/Q _14215_/Q _14151_/Q _14469_/Q _12641_/S _12689_/S1 vssd1 vssd1
+ vccd1 vccd1 _12639_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _15427_/CLK hold918/X vssd1 vssd1 vccd1 vccd1 hold917/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11697__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14309_ _15268_/CLK hold818/X vssd1 vssd1 vccd1 vccd1 hold817/A sky130_fd_sc_hd__dfxtp_1
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13478__A _13487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15289_ _15289_/CLK hold964/X vssd1 vssd1 vccd1 vccd1 hold963/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08071__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__B _13197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09003__A2 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09634__S0 _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07014__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2522_A _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _10002_/C _10110_/A _10283_/C _10115_/D vssd1 vssd1 vccd1 vccd1 _09851_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__08211__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10106__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout707 hold465/X vssd1 vssd1 vccd1 vccd1 _13690_/A1 sky130_fd_sc_hd__buf_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 _12329_/A vssd1 vssd1 vccd1 vccd1 _13651_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout729 _14959_/Q vssd1 vssd1 vccd1 vccd1 _10283_/C sky130_fd_sc_hd__buf_6
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__and2b_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _13665_/A1 hold1329/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06993_/X sky130_fd_sc_hd__mux2_1
X_09781_ _10233_/A _09923_/B _09781_/C vssd1 vssd1 vccd1 vccd1 _09781_/X sky130_fd_sc_hd__or3_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08732_ _08630_/A _08628_/A _08629_/A vssd1 vssd1 vccd1 vccd1 _08734_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11649__A1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ hold803/A _14537_/Q _14697_/Q _14761_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08663_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07614_ hold1831/X _13687_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07614_/X sky130_fd_sc_hd__mux2_1
X_08594_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08597_/A sky130_fd_sc_hd__xor2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07545_ _13386_/A hold173/X vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_127_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15446_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout438_A _07644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10624__A2 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07476_ _14088_/Q _14089_/Q _11729_/C vssd1 vssd1 vccd1 vccd1 _07778_/B sky130_fd_sc_hd__or3_4
XFILLER_0_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12276__B _12276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09215_ _09215_/A _09215_/B vssd1 vssd1 vccd1 vccd1 _09217_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_173_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10077__A _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout605_A _15209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _09146_/A _09146_/B _09146_/C vssd1 vssd1 vccd1 vccd1 _09317_/A sky130_fd_sc_hd__or3_2
XANTENNA__09866__A _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13388__A _13393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _12221_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12129__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08028_ _07965_/Y _08024_/X _08027_/Y vssd1 vssd1 vccd1 vccd1 _08028_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_124_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold750 hold750/A vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 hold761/A vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 hold772/A vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold783 hold783/A vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 hold794/A vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ _10183_/A _09979_/B _09979_/C _09979_/D vssd1 vssd1 vccd1 vccd1 _10182_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2140 _07756_/X vssd1 vssd1 vccd1 vccd1 _14372_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2151 _13800_/Q vssd1 vssd1 vccd1 vccd1 hold2151/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2162 _13503_/X vssd1 vssd1 vccd1 vccd1 _15261_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2173 _14457_/Q vssd1 vssd1 vccd1 vccd1 hold2173/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ hold309/X hold759/X _12991_/S vssd1 vssd1 vccd1 vccd1 _12990_/X sky130_fd_sc_hd__mux2_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2184 _07132_/X vssd1 vssd1 vccd1 vccd1 _13942_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07939__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1450 _07693_/X vssd1 vssd1 vccd1 vccd1 _14313_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2195 _14529_/Q vssd1 vssd1 vccd1 vccd1 hold2195/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1461 _14545_/Q vssd1 vssd1 vccd1 vccd1 hold1461/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _13729_/A1 hold1961/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11941_/X sky130_fd_sc_hd__mux2_1
Xhold1472 _11970_/X vssd1 vssd1 vccd1 vccd1 _14789_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1483 _14514_/Q vssd1 vssd1 vccd1 vccd1 hold1483/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 _11802_/X vssd1 vssd1 vccd1 vccd1 _14626_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14660_ _15042_/CLK _14660_/D vssd1 vssd1 vccd1 vccd1 _14660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ hold579/X _13693_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold580/A sky130_fd_sc_hd__mux2_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ input62/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__or2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _11378_/D _10822_/X _10821_/X vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__13570__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__A2 _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15374_/CLK sky130_fd_sc_hd__clkbuf_16
X_14591_ _15390_/CLK _14591_/D vssd1 vssd1 vccd1 vccd1 _14591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_211_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10076__B1 _07319_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _14427_/Q _13590_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
XFILLER_0_165_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ _15159_/Q _07812_/A _13590_/B _10753_/X vssd1 vssd1 vccd1 vccd1 _10754_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07060__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _10684_/A _10684_/B _10684_/C vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13473_ _13481_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__and2_2
XFILLER_0_192_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08116__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__B1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15212_ _15429_/CLK _15212_/D vssd1 vssd1 vccd1 vccd1 _15212_/Q sky130_fd_sc_hd__dfxtp_1
X_12424_ _13866_/Q _13994_/Q hold809/A hold929/A _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12424_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15143_ _15304_/CLK _15143_/D vssd1 vssd1 vccd1 vccd1 _15143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _12379_/A _12379_/B _13375_/B vssd1 vssd1 vccd1 vccd1 _12355_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08992__A1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11306_ _14811_/Q hold875/A hold341/A _14747_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _11307_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15074_ _15432_/CLK _15074_/D vssd1 vssd1 vccd1 vccd1 _15074_/Q sky130_fd_sc_hd__dfxtp_1
X_12286_ _13455_/A _12286_/B vssd1 vssd1 vccd1 vccd1 _14935_/D sky130_fd_sc_hd__and2_2
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11237_ _11567_/A _15226_/Q vssd1 vssd1 vccd1 vccd1 _11239_/B sky130_fd_sc_hd__nand2_1
X_14025_ _15351_/CLK hold314/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11168_ _11168_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_184_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10119_ _10119_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__xnor2_2
X_11099_ _11281_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10450__A _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12828__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12923__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ _15247_/CLK _14927_/D vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11980__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14858_ _15004_/CLK _14858_/D vssd1 vssd1 vccd1 vccd1 _14858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13809_ _15080_/CLK _13809_/D vssd1 vssd1 vccd1 vccd1 _13809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_109_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15379_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ _15079_/CLK _14789_/D vssd1 vssd1 vccd1 vccd1 _14789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08574__B _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07330_ _08102_/A _07330_/B _07330_/C _07330_/D vssd1 vssd1 vccd1 vccd1 _07330_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__08355__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07261_ _07261_/A _07261_/B vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09000_ _09726_/B _09124_/B vssd1 vssd1 vccd1 vccd1 _09127_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13700__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__S0 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07192_ hold1705/X _13512_/A0 _07198_/S vssd1 vssd1 vccd1 vccd1 _07192_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_171_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2737_A _15189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07918__B _07919_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13001__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09902_ _09747_/X _09749_/Y _09900_/Y _09901_/X vssd1 vssd1 vccd1 vccd1 _09903_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout504 _13092_/A1 vssd1 vssd1 vccd1 vccd1 _12917_/A1 sky130_fd_sc_hd__buf_6
Xfanout515 _11497_/A vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout526 _11499_/B1 vssd1 vssd1 vccd1 vccd1 _11510_/A1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07934__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09833_ _09833_/A _09833_/B _09833_/C vssd1 vssd1 vccd1 vccd1 _09833_/X sky130_fd_sc_hd__and3_2
Xfanout537 _15424_/Q vssd1 vssd1 vccd1 vccd1 _11507_/A sky130_fd_sc_hd__buf_6
Xfanout548 _10425_/S1 vssd1 vssd1 vccd1 vccd1 _10087_/S1 sky130_fd_sc_hd__buf_6
Xfanout559 _08763_/S0 vssd1 vssd1 vccd1 vccd1 _08990_/S0 sky130_fd_sc_hd__buf_8
XANTENNA_fanout388_A _11696_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09764_/X sky130_fd_sc_hd__or2_1
X_06976_ _07875_/B _07114_/B vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07145__S _07147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08715_ _08714_/B _08714_/C _08714_/A vssd1 vssd1 vccd1 vccd1 _08717_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__12914__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09695_ _09555_/B _09557_/B _09693_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _09745_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout555_A _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__A0 _13705_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ _13558_/A _09222_/B hold2533/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _14435_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13390__B _13390_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14917__D _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ _08901_/A _09866_/B _08577_/C vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__and3_1
XFILLER_0_117_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout722_A _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11191__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09999__B1 _14963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07528_ hold605/X _13732_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 hold606/A sky130_fd_sc_hd__mux2_1
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ _07459_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14089_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08671__B1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ _11537_/B _10468_/X _10469_/X vssd1 vssd1 vccd1 vccd1 _10472_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08649__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ _09271_/A _09129_/B vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__or2_1
XFILLER_0_161_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _14881_/Q _12172_/B vssd1 vssd1 vccd1 vccd1 _12140_/X sky130_fd_sc_hd__or2_1
XANTENNA__08974__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ hold2481/X _12099_/A2 _12070_/X _13492_/A vssd1 vssd1 vccd1 vccd1 _12071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 hold580/A vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 hold591/A vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _11022_/A _11022_/B _11022_/C vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07055__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ hold241/A hold961/A hold1245/X _13984_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12973_/X sky130_fd_sc_hd__mux4_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1280 _07777_/X vssd1 vssd1 vccd1 vccd1 _14393_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1291 _14399_/Q vssd1 vssd1 vccd1 vccd1 hold1291/X sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ _14776_/CLK _14712_/D vssd1 vssd1 vccd1 vccd1 _14712_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _13679_/A1 hold2009/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11924_/X sky130_fd_sc_hd__mux2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _15372_/CLK _14643_/D vssd1 vssd1 vccd1 vccd1 _14643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ hold1077/X _13742_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10806_ _11573_/A _11605_/B _10807_/C _10807_/D vssd1 vssd1 vccd1 vccd1 _10806_/Y
+ sky130_fd_sc_hd__a22oi_2
X_14574_ _15373_/CLK hold224/X vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11786_ hold507/X _13673_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold508/A sky130_fd_sc_hd__mux2_1
XFILLER_0_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12994__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13525_ _13673_/A1 hold951/X _13534_/S vssd1 vssd1 vccd1 vccd1 hold952/A sky130_fd_sc_hd__mux2_1
X_10737_ _10395_/B _10736_/Y _10735_/Y vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13520__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _13468_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _13456_/Y sky130_fd_sc_hd__nand2_1
X_10668_ _10668_/A _10668_/B _10464_/B vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _12482_/A _12407_/B vssd1 vssd1 vccd1 vccd1 _14944_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _07274_/B _07280_/B _07274_/A vssd1 vssd1 vccd1 vccd1 _10599_/X sky130_fd_sc_hd__a21bo_1
X_13387_ _13393_/A _13387_/B vssd1 vssd1 vccd1 vccd1 _15178_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10221__B1 _11474_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__A1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15126_ _15132_/CLK _15126_/D vssd1 vssd1 vccd1 vccd1 _15126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _15391_/Q _14526_/Q hold343/A _14750_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12338_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11975__S _11977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _15190_/CLK _15057_/D vssd1 vssd1 vccd1 vccd1 _15057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ _13168_/A _13424_/B vssd1 vssd1 vccd1 vccd1 _14918_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14008_ _15087_/CLK _14008_/D vssd1 vssd1 vccd1 vccd1 _14008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07473__B _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08500_ _08500_/A _08500_/B _08500_/C vssd1 vssd1 vccd1 vccd1 _08502_/A sky130_fd_sc_hd__and3_1
XFILLER_0_204_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09480_ _07243_/B _09340_/A _09340_/B _07241_/Y vssd1 vssd1 vccd1 vccd1 _09481_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08585__A _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08431_ _08378_/X _08379_/Y _08430_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _13383_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _12247_/A _08359_/X _08361_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _08363_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ _09437_/A _11351_/B vssd1 vssd1 vccd1 vccd1 _07313_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08293_ _09008_/A _08809_/B _08809_/D _08893_/A vssd1 vssd1 vccd1 vccd1 _08294_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07244_ _09864_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _09133_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_160_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07208__A1 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07175_ _11921_/A0 hold1873/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07175_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12201__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__A0 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11885__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09863__B _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13385__B _13385_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__C _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _09816_/A _10338_/C vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__nand2_1
Xfanout367 _12259_/A1 vssd1 vssd1 vccd1 vccd1 _11514_/B1 sky130_fd_sc_hd__buf_8
Xfanout378 _12323_/X vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__clkbuf_16
Xfanout389 _11652_/Y vssd1 vssd1 vccd1 vccd1 _11668_/S sky130_fd_sc_hd__clkbuf_16
X_09747_ _09601_/C _09602_/X _09744_/Y _09746_/X vssd1 vssd1 vccd1 vccd1 _09747_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06959_ _07453_/A _06950_/B _06958_/X _06953_/X vssd1 vssd1 vccd1 vccd1 _06959_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12363__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08495__A _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _10185_/A _09979_/C _09678_/C _09824_/A vssd1 vssd1 vccd1 vccd1 _09824_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07603__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08629_/A _08629_/B vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__nand2_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ hold2784/X _11283_/S _11640_/B1 vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__o21a_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11243__A2 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11571_ _11441_/A _11441_/B _11441_/C _11445_/C vssd1 vssd1 vccd1 vccd1 _11572_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ input79/X fanout2/X _13309_/X vssd1 vssd1 vccd1 vccd1 _13311_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10522_ _10522_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__xor2_2
X_14290_ _15451_/CLK hold426/X vssd1 vssd1 vccd1 vccd1 hold425/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10453_ _11597_/A _11605_/B _10277_/B _10275_/X vssd1 vssd1 vccd1 vccd1 _10455_/B
+ sky130_fd_sc_hd__a31o_1
X_13241_ _13241_/A _13241_/B _13241_/C _13241_/D vssd1 vssd1 vccd1 vccd1 fanout4/A
+ sky130_fd_sc_hd__and4_4
XFILLER_0_134_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10429__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10384_ _10201_/X _10204_/Y _10382_/Y _10383_/X vssd1 vssd1 vccd1 vccd1 _10387_/A
+ sky130_fd_sc_hd__a211oi_2
X_13172_ _13178_/A _13172_/B vssd1 vssd1 vccd1 vccd1 _15037_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11795__S _11795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ hold2489/X _12129_/A2 _12122_/X _12063_/A vssd1 vssd1 vccd1 vccd1 _12123_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _12120_/A hold2699/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07574__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _11536_/A _11623_/A _11537_/B _11542_/A vssd1 vssd1 vccd1 vccd1 _11010_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout890 _13317_/A vssd1 vssd1 vccd1 vccd1 _12482_/A sky130_fd_sc_hd__buf_4
XANTENNA__12259__A1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__B2 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08558__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ _13106_/A1 _13165_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12957_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09675__A2 _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07513__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _13662_/A1 hold2263/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__mux2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12887_ _13024_/S1 _12884_/X _12886_/X vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__a21o_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _15042_/CLK _14626_/D vssd1 vssd1 vccd1 vccd1 _14626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ hold1787/X _13725_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/CLK hold166/X vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12431__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ hold1341/X _13656_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15222_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _13689_/A1 hold2121/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13508_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _15348_/CLK _14488_/D vssd1 vssd1 vccd1 vccd1 _14488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_183_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12719__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ _09213_/B _13440_/S _13438_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15213_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09386__D _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10606__C _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15116_/CLK _15109_/D vssd1 vssd1 vccd1 vccd1 _15109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13486__A _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ hold937/A hold669/A _14636_/Q _14732_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08981_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2706 _15127_/Q vssd1 vssd1 vccd1 vccd1 hold2706/X sky130_fd_sc_hd__dlygate4sd3_1
X_07931_ _08197_/A _07928_/X _07930_/X vssd1 vssd1 vccd1 vccd1 _07931_/Y sky130_fd_sc_hd__o21ai_1
Xhold2717 _12052_/X vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2728 _15058_/Q vssd1 vssd1 vccd1 vccd1 hold2728/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2739 _15180_/Q vssd1 vssd1 vccd1 vccd1 hold2739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07862_ _07862_/A _07862_/B _07862_/C _07862_/D vssd1 vssd1 vccd1 vccd1 _07862_/X
+ sky130_fd_sc_hd__and4_4
XANTENNA__11170__A1 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09601_ _09602_/A _09602_/B _09601_/C _09601_/D vssd1 vssd1 vccd1 vccd1 _09601_/X
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__11170__B2 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07793_ hold1833/X _13698_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 _07793_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09115__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09204__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09464_/A _09464_/B _09464_/C vssd1 vssd1 vccd1 vccd1 _09463_/X sky130_fd_sc_hd__and3_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ _08474_/A _08413_/C _08413_/A vssd1 vssd1 vccd1 vccd1 _08415_/C sky130_fd_sc_hd__a21o_1
X_09394_ _09395_/A _09395_/B vssd1 vssd1 vccd1 vccd1 _09394_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_191_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09858__B _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A _13650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15392_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout518_A _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ _08873_/A _08276_/B vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12284__B _12284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10984__A1 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10984__B2 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07227_ _08496_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _08102_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ _13725_/A1 hold1749/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07158_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout887_A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13396__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14930__D _14930_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ _13725_/A1 hold2287/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07089_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_98_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _14987_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09354__A1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12810_ _14673_/Q _13946_/Q _12841_/S vssd1 vssd1 vccd1 vccd1 _12810_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12336__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13790_ _06905_/A _13792_/A2 _11689_/X _07450_/B vssd1 vssd1 vccd1 vccd1 _15348_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09114__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _14347_/Q _14251_/Q _12741_/S vssd1 vssd1 vccd1 vccd1 _12741_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ _15460_/CLK _15460_/D vssd1 vssd1 vccd1 vccd1 _15460_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12672_ hold639/A _14507_/Q hold887/A _14731_/Q _12641_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12672_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_182_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14411_ _15375_/CLK hold978/X vssd1 vssd1 vccd1 vccd1 hold977/A sky130_fd_sc_hd__dfxtp_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11623_ _11623_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11624_/S sky130_fd_sc_hd__nand2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12413__A1 _12642_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ _15391_/CLK _15391_/D vssd1 vssd1 vccd1 vccd1 _15391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15261_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_167_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07569__A _13396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14342_ _15372_/CLK _14342_/D vssd1 vssd1 vccd1 vccd1 _14342_/Q sky130_fd_sc_hd__dfxtp_1
X_11554_ _11554_/A _11554_/B vssd1 vssd1 vccd1 vccd1 _11555_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10505_ _10295_/Y _10332_/X _10502_/Y _10503_/X vssd1 vssd1 vccd1 vccd1 _10505_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07288__B _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14273_ _15080_/CLK _14273_/D vssd1 vssd1 vccd1 vccd1 _14273_/Q sky130_fd_sc_hd__dfxtp_1
X_11485_ _13750_/A _13372_/B vssd1 vssd1 vccd1 vccd1 _11485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ hold1017/X _13736_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 _13224_/X sky130_fd_sc_hd__mux2_1
X_10436_ _07280_/B _10262_/X _10600_/A vssd1 vssd1 vccd1 vccd1 _10436_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_output172_A _15184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08396__A2 _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13155_ _13389_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _15020_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_209_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10367_ _10189_/B _10191_/B _10364_/X _10365_/Y vssd1 vssd1 vccd1 vccd1 _10367_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12106_ _14993_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12106_/X
+ sky130_fd_sc_hd__or4_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07508__S _07509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10298_ _11614_/A _10827_/C _10827_/D _11586_/A vssd1 vssd1 vccd1 vccd1 _10298_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13086_ _13092_/A1 _13085_/X _13100_/S0 vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10442__B _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15389_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12037_ _12037_/A _12037_/B vssd1 vssd1 vccd1 vccd1 _14831_/D sky130_fd_sc_hd__and2_1
XANTENNA__12575__S1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11152__A1 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__B2 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _15384_/CLK _13988_/D vssd1 vssd1 vccd1 vccd1 _13988_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09024__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _14291_/Q _14227_/Q hold477/A _14481_/Q _12915_/S _12939_/S1 vssd1 vssd1
+ vccd1 vccd1 _12939_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_158_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14609_ _15376_/CLK _14609_/D vssd1 vssd1 vccd1 vccd1 _14609_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09678__B _09979_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12404__A1 _13377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2385_A _14429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08582__B _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15460_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ hold641/A _14531_/Q _14691_/Q _14755_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _08130_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08084__A1 _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10966__A1 _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10617__B _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__B2 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ _08981_/A _08061_/B vssd1 vssd1 vccd1 vccd1 _08061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2552_A _14453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07012_ _07182_/A _13716_/A vssd1 vssd1 vccd1 vccd1 _07012_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_4_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__A1 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _11288_/A1 _13388_/B _08884_/X vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__a21oi_4
Xhold2503 _10085_/X vssd1 vssd1 vccd1 vccd1 _14446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2514 _12073_/X vssd1 vssd1 vccd1 vccd1 _14848_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09336__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2525 _15353_/Q vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07914_ _07908_/B _07908_/C _07908_/A vssd1 vssd1 vccd1 vccd1 _07915_/B sky130_fd_sc_hd__a21o_1
Xhold2536 _12185_/X vssd1 vssd1 vccd1 vccd1 _14903_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1802 _06997_/X vssd1 vssd1 vccd1 vccd1 _13816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2547 _15033_/Q vssd1 vssd1 vccd1 vccd1 _07573_/B sky130_fd_sc_hd__dlygate4sd3_1
X_08894_ _09136_/A _09866_/B _08895_/C _08895_/D vssd1 vssd1 vccd1 vccd1 _08894_/X
+ sky130_fd_sc_hd__and4_1
Xhold1813 _15411_/Q vssd1 vssd1 vccd1 vccd1 hold1813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2558 _15117_/Q vssd1 vssd1 vccd1 vccd1 hold2558/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10577__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2569 hold2859/X vssd1 vssd1 vccd1 vccd1 hold2569/X sky130_fd_sc_hd__buf_1
Xhold1824 _07057_/X vssd1 vssd1 vccd1 vccd1 _13873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1835 _14247_/Q vssd1 vssd1 vccd1 vccd1 hold1835/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ _07862_/B _14032_/Q _07841_/X _07843_/X _07844_/X vssd1 vssd1 vccd1 vccd1
+ _07846_/C sky130_fd_sc_hd__o2111a_1
Xhold1846 _13515_/X vssd1 vssd1 vccd1 vccd1 _15273_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11694__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1857 _14805_/Q vssd1 vssd1 vccd1 vccd1 hold1857/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout370_A _07899_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1868 _13669_/X vssd1 vssd1 vccd1 vccd1 _15376_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout468_A _07884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1879 _13842_/Q vssd1 vssd1 vccd1 vccd1 hold1879/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12318__S1 _12343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07776_ _13681_/A1 hold1129/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07776_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07153__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__B _13444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ hold879/A _14544_/Q _14704_/Q _14768_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09515_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_196_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12643__A1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ _10115_/A _09726_/B _09445_/C _09579_/A vssd1 vssd1 vccd1 vccd1 _09447_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06992__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _11320_/A _09377_/B vssd1 vssd1 vccd1 vccd1 _09377_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout802_A _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14925__D _14925_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ _08420_/A _08327_/B _08327_/C vssd1 vssd1 vccd1 vccd1 _08329_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08259_ _14430_/Q _13546_/A _08049_/B _08257_/A vssd1 vssd1 vccd1 vccd1 _08259_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11270_ _11465_/A _11269_/B _11269_/C vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_104_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ _10219_/Y _10220_/X _11474_/A2 vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__a21o_1
X_10152_ _10152_/A _10152_/B _10152_/C vssd1 vssd1 vccd1 vccd1 _10154_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09109__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput290 _14885_/Q vssd1 vssd1 vccd1 vccd1 out0[8] sky130_fd_sc_hd__buf_12
X_14960_ _14971_/CLK _14960_/D vssd1 vssd1 vccd1 vccd1 _14960_/Q sky130_fd_sc_hd__dfxtp_1
X_10083_ _13580_/A _10082_/B _10232_/B _10233_/A vssd1 vssd1 vccd1 vccd1 _10083_/Y
+ sky130_fd_sc_hd__a211oi_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ _15444_/CLK _13911_/D vssd1 vssd1 vccd1 vccd1 _13911_/Q sky130_fd_sc_hd__dfxtp_1
X_14891_ _14989_/CLK _14891_/D vssd1 vssd1 vccd1 vccd1 _14891_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13065__S _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07984__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ _14569_/CLK _13842_/D vssd1 vssd1 vccd1 vccd1 _13842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ hold223/X vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10985_ _11590_/A _11573_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _10987_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_70_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08302__A2 _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12724_ _13878_/Q _14006_/Q _13846_/Q _13814_/Q _12791_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12724_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08683__A _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _15443_/CLK hold396/X vssd1 vssd1 vccd1 vccd1 hold395/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ _12327_/A _12654_/X _12652_/X vssd1 vssd1 vccd1 vccd1 _13153_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12409__S _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11606_ _11606_/A _11606_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13595__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15374_ _15374_/CLK hold768/X vssd1 vssd1 vccd1 vccd1 hold767/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12586_ _12642_/A1 _12585_/X _12700_/S0 vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14325_ _14926_/CLK _14325_/D vssd1 vssd1 vccd1 vccd1 _14325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11537_ _11537_/A _11537_/B vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold409 hold409/A vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14256_ _15062_/CLK hold700/X vssd1 vssd1 vccd1 vccd1 hold699/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11468_ _11468_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__or2_1
XFILLER_0_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__A1 _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ hold2111/X _13653_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13207_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09566__B2 _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ hold299/A hold431/A hold295/A _14742_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10420_/B sky130_fd_sc_hd__mux4_1
X_14187_ _15278_/CLK hold120/X vssd1 vssd1 vccd1 vccd1 _14187_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12796__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10176__A2 _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _11399_/A _11399_/B _11399_/C vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__and3_1
XFILLER_0_21_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13499_/A hold171/X vssd1 vssd1 vccd1 vccd1 hold172/A sky130_fd_sc_hd__and2_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11983__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12548__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13100_/S0 _13064_/X _13068_/X _13100_/S1 vssd1 vssd1 vccd1 vccd1 _13070_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15433_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1109 _14342_/Q vssd1 vssd1 vccd1 vccd1 hold1109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold2300_A _13473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ hold1433/X _13736_/A1 _07642_/S vssd1 vssd1 vccd1 vccd1 _07630_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07561_ _13396_/A hold177/X vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__and2_1
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09300_ _09542_/A _11561_/A _10022_/B _09858_/C vssd1 vssd1 vccd1 vccd1 _09400_/A
+ sky130_fd_sc_hd__nand4_4
XANTENNA__13703__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07492_ hold1811/X _13698_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07492_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07701__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ _09514_/A _09228_/X _09230_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09232_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12928__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ _09162_/A _09162_/B vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ _13546_/A _08441_/B hold2640/X _13178_/A vssd1 vssd1 vccd1 vccd1 _14429_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09093_ _09087_/A _09222_/B _09092_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _09093_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08044_ _14427_/Q _14426_/Q _14428_/Q vssd1 vssd1 vccd1 vccd1 _08044_/X sky130_fd_sc_hd__a21o_1
Xhold910 hold910/A vssd1 vssd1 vccd1 vccd1 hold910/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold921 hold921/A vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 hold932/A vssd1 vssd1 vccd1 vccd1 hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 hold943/A vssd1 vssd1 vccd1 vccd1 hold943/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 hold954/A vssd1 vssd1 vccd1 vccd1 hold954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 hold965/A vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__B1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 hold976/A vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold987 hold987/A vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 hold998/A vssd1 vssd1 vccd1 vccd1 hold998/X sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _09995_/A _09995_/B _09995_/C vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__or3_2
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout585_A _10166_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__C1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2300 _13473_/X vssd1 vssd1 vccd1 vccd1 _15232_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2311 _15015_/Q vssd1 vssd1 vccd1 vccd1 _07555_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11893__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2322 _14997_/Q vssd1 vssd1 vccd1 vccd1 _12114_/A sky130_fd_sc_hd__buf_2
XFILLER_0_196_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08946_ _08829_/B _08829_/Y _08944_/Y _08945_/X vssd1 vssd1 vccd1 vccd1 _08948_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12539__S1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2333 hold2851/X vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06987__S _06994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__A1 _10233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2344 _13545_/X vssd1 vssd1 vccd1 vccd1 _15298_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2355 _13339_/Y vssd1 vssd1 vccd1 vccd1 _13340_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1610 _13530_/X vssd1 vssd1 vccd1 vccd1 _15288_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2366 _13751_/X vssd1 vssd1 vccd1 vccd1 hold2366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 _14228_/Q vssd1 vssd1 vccd1 vccd1 hold1621/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13393__B _13393_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1632 _11657_/X vssd1 vssd1 vccd1 vccd1 _14460_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2377 _07949_/X vssd1 vssd1 vccd1 vccd1 hold2377/X sky130_fd_sc_hd__dlygate4sd3_1
X_08877_ _08877_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _08877_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout752_A _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2388 _15324_/Q vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__buf_1
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1643 _15394_/Q vssd1 vssd1 vccd1 vccd1 hold1643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2399 _12097_/X vssd1 vssd1 vccd1 vccd1 _14860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1654 _07047_/X vssd1 vssd1 vccd1 vccd1 _13863_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1665 _14213_/Q vssd1 vssd1 vccd1 vccd1 hold1665/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _08873_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07828_/Y sky130_fd_sc_hd__nor2_1
Xhold1676 _07728_/X vssd1 vssd1 vccd1 vccd1 _14347_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1687 _13857_/Q vssd1 vssd1 vccd1 vccd1 hold1687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1698 _11808_/X vssd1 vssd1 vccd1 vccd1 _14632_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07759_ _13664_/A1 hold1593/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _14680_/Q _13953_/Q hold715/A _13921_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10771_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07611__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09429_ _10022_/A _14950_/Q _09858_/B _10142_/B vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12440_ hold1291/X hold1113/X _12441_/S vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09245__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12475__S0 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _15360_/Q _15263_/Q _15071_/Q _14364_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12371_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ _15434_/CLK _14110_/D vssd1 vssd1 vccd1 vccd1 _14110_/Q sky130_fd_sc_hd__dfxtp_1
X_11322_ _13714_/A1 _07899_/Y _07900_/Y _13202_/B _11320_/Y vssd1 vssd1 vccd1 vccd1
+ _11322_/X sky130_fd_sc_hd__a221o_1
X_15090_ _15090_/CLK _15090_/D vssd1 vssd1 vccd1 vccd1 _15090_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13568__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14041_ _14042_/CLK _14041_/D vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
X_11253_ _11252_/B _11252_/C _11252_/A vssd1 vssd1 vccd1 vccd1 _11254_/C sky130_fd_sc_hd__a21o_1
XANTENNA__10273__A _14964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07058__S _07061_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _10206_/C vssd1 vssd1 vccd1 vccd1 _10204_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11184_ _11183_/A _11183_/B _11371_/B _11183_/D vssd1 vssd1 vccd1 vccd1 _11184_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _10306_/A _11168_/A _10135_/C _10135_/D vssd1 vssd1 vccd1 vccd1 _10135_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_24_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10066_ _10065_/B _10065_/C _10065_/A vssd1 vssd1 vccd1 vccd1 _10066_/Y sky130_fd_sc_hd__a21oi_1
X_14943_ _15392_/CLK _14943_/D vssd1 vssd1 vccd1 vccd1 _14943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12855__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ _14876_/CLK _14874_/D vssd1 vssd1 vccd1 vccd1 _14874_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12950__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13825_ _15385_/CLK _13825_/D vssd1 vssd1 vccd1 vccd1 _13825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13523__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13756_ hold165/X vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__clkbuf_1
X_10968_ _11598_/A _11594_/B _10969_/C _11150_/A vssd1 vssd1 vccd1 vccd1 _10970_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06926__A _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__B2 _13180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12707_ _13150_/A _12707_/B vssd1 vssd1 vccd1 vccd1 _14956_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_39_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10448__A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ hold1333/X _13687_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 _13687_/X sky130_fd_sc_hd__mux2_1
X_10899_ _10896_/A _10897_/X _10713_/B _10713_/Y vssd1 vssd1 vccd1 vccd1 _10900_/D
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__09659__D _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15426_ _15426_/CLK _15426_/D vssd1 vssd1 vccd1 vccd1 _15426_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12638_ _12642_/B1 _12633_/X _12637_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12645_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11978__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15357_ _15357_/CLK _15357_/D vssd1 vssd1 vccd1 vccd1 _15357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12240__C1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _12669_/A1 _12564_/X _12568_/X _12700_/S1 vssd1 vssd1 vccd1 vccd1 _12570_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14308_ _15400_/CLK hold506/X vssd1 vssd1 vccd1 vccd1 hold505/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ _15385_/CLK _15288_/D vssd1 vssd1 vccd1 vccd1 _15288_/Q sky130_fd_sc_hd__dfxtp_1
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ _15391_/CLK _14239_/D vssd1 vssd1 vccd1 vccd1 _14239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10183__A _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09634__S1 _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09972__A _14941_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__A1 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08211__B2 _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 _13689_/A1 vssd1 vssd1 vccd1 vccd1 _13656_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout719 hold2415/X vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__buf_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08800_/A _08800_/B vssd1 vssd1 vccd1 vccd1 _08802_/B sky130_fd_sc_hd__xnor2_2
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13494__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09780_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09781_/C sky130_fd_sc_hd__nor2_1
X_06992_ _13664_/A1 hold1315/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06992_/X sky130_fd_sc_hd__mux2_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08841_/A _08731_/B vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__and2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08662_ _08989_/A _08662_/B vssd1 vssd1 vccd1 vccd1 _08662_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ hold327/X _13719_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 hold328/A sky130_fd_sc_hd__mux2_1
XFILLER_0_205_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08593_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08593_/X sky130_fd_sc_hd__and2_1
XFILLER_0_178_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07544_ hold1235/X _13715_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 _07544_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07475_ hold65/X _07475_/B vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__and2_1
XFILLER_0_119_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10358__A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13559__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09214_ _09213_/B _09214_/B vssd1 vssd1 vccd1 vccd1 _09215_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11888__S _11893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ _09145_/A _09145_/B vssd1 vssd1 vccd1 vccd1 _09146_/C sky130_fd_sc_hd__and2_1
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout500_A _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09076_ _09075_/A _09075_/C _09075_/B vssd1 vssd1 vccd1 vccd1 _09205_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13388__B _13388_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12209__S0 _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08027_ _07965_/Y _08024_/X _10397_/A vssd1 vssd1 vccd1 vccd1 _08027_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11189__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold740 hold740/A vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 hold751/A vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold762 hold762/A vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap481 _07359_/B vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__clkbuf_2
Xhold773 hold773/A vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold784 hold784/A vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 hold795/A vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ _09979_/B _09979_/C _09979_/D _10183_/A vssd1 vssd1 vccd1 vccd1 _09981_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2130 _11919_/X vssd1 vssd1 vccd1 vccd1 _14740_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2141 _14363_/Q vssd1 vssd1 vccd1 vccd1 hold2141/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07606__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08929_ _09039_/B _08928_/C _08928_/A vssd1 vssd1 vccd1 vccd1 _08930_/C sky130_fd_sc_hd__a21o_1
Xhold2152 _06981_/X vssd1 vssd1 vccd1 vccd1 _13800_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2163 _14528_/Q vssd1 vssd1 vccd1 vccd1 hold2163/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12837__A1 _12939_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2174 _11654_/X vssd1 vssd1 vccd1 vccd1 _14457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1440 _11950_/X vssd1 vssd1 vccd1 vccd1 _14770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2185 _13916_/Q vssd1 vssd1 vccd1 vccd1 hold2185/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 _14019_/Q vssd1 vssd1 vccd1 vccd1 hold1451/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _13728_/A1 hold2127/X _11943_/S vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__mux2_1
Xhold2196 _11735_/X vssd1 vssd1 vccd1 vccd1 _14529_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1462 _11751_/X vssd1 vssd1 vccd1 vccd1 _14545_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1473 _15074_/Q vssd1 vssd1 vccd1 vccd1 hold1473/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1484 _11718_/X vssd1 vssd1 vccd1 vccd1 _14514_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1495 _13819_/Q vssd1 vssd1 vccd1 vccd1 hold1495/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ hold815/X _13725_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold816/A sky130_fd_sc_hd__mux2_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13610_ _07428_/A _13625_/C _13609_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _15332_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10822_ _11586_/A _11614_/A _11378_/C vssd1 vssd1 vccd1 vccd1 _10822_/X sky130_fd_sc_hd__and3_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08269__A1 _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13262__A1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _15299_/CLK hold908/X vssd1 vssd1 vccd1 vccd1 hold907/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12696__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08364__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _15296_/D sky130_fd_sc_hd__and2_1
XFILLER_0_177_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10753_ _13588_/A _10751_/B _10752_/Y _07390_/A vssd1 vssd1 vccd1 vccd1 _10753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_165_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _13481_/A _13472_/B vssd1 vssd1 vccd1 vccd1 _13472_/X sky130_fd_sc_hd__and2_1
XFILLER_0_165_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10684_ _10684_/A _10684_/B _10684_/C vssd1 vssd1 vccd1 vccd1 _10686_/A sky130_fd_sc_hd__and3_1
XANTENNA__12448__S0 _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11798__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15211_ _15429_/CLK _15211_/D vssd1 vssd1 vccd1 vccd1 _15211_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09769__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ hold185/A _14302_/Q hold861/A _13962_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12423_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08116__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12999__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11120__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15142_ _15301_/CLK _15142_/D vssd1 vssd1 vccd1 vccd1 _15142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ _12326_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12354_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ hold953/A hold677/A hold451/A _14392_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _11305_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15073_ _15265_/CLK _15073_/D vssd1 vssd1 vccd1 vccd1 _15073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _13171_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _14934_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_121_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14024_ _15348_/CLK hold282/X vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09792__A _10244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _11236_/A _11236_/B vssd1 vssd1 vccd1 vccd1 _11239_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_205_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13518__S _13518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11167_ _11606_/B _11166_/X _11165_/X vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07952__B1 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07516__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ _11590_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11098_ _11098_/A _11098_/B _11096_/Y vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__or3b_1
XANTENNA__10450__B _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10839__B1 _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10049_ _10046_/X _10047_/Y _09885_/Y _09887_/X vssd1 vssd1 vccd1 vccd1 _10050_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12923__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08052__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14926_ _14926_/CLK _14926_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11500__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10934__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14857_ _15004_/CLK _14857_/D vssd1 vssd1 vccd1 vccd1 _14857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13808_ _15079_/CLK _13808_/D vssd1 vssd1 vccd1 vccd1 _13808_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13253__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14788_ _15365_/CLK _14788_/D vssd1 vssd1 vccd1 vccd1 _14788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08574__C _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13739_ hold1947/X _13739_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 _13739_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08355__S1 _12244_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09967__A _14942_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ _11614_/B _10108_/C vssd1 vssd1 vccd1 vccd1 _07261_/B sky130_fd_sc_hd__or2_1
XANTENNA__13005__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12439__S0 _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08871__A _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11016__B1 _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15409_ _15446_/CLK hold880/X vssd1 vssd1 vccd1 vccd1 hold879/A sky130_fd_sc_hd__dfxtp_1
X_07191_ hold421/X _13659_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold422/A sky130_fd_sc_hd__mux2_1
XANTENNA__13100__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_83_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08432__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10775__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2632_A _15460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ _09898_/Y _09899_/X _09693_/Y _09696_/Y vssd1 vssd1 vccd1 vccd1 _09901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _06942_/Y vssd1 vssd1 vccd1 vccd1 _13092_/A1 sky130_fd_sc_hd__buf_6
Xfanout516 _10252_/A vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__buf_6
X_09832_ _09831_/B _09831_/C _09831_/A vssd1 vssd1 vccd1 vccd1 _09833_/C sky130_fd_sc_hd__a21o_1
Xfanout527 _10255_/A1 vssd1 vssd1 vccd1 vccd1 _11499_/B1 sky130_fd_sc_hd__buf_4
Xfanout538 _08763_/S1 vssd1 vssd1 vccd1 vccd1 _08548_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_141_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _10425_/S1 vssd1 vssd1 vccd1 vccd1 _09795_/S1 sky130_fd_sc_hd__clkbuf_8
X_09763_ _09763_/A _09763_/B vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12819__A1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ _07875_/C _07643_/C vssd1 vssd1 vccd1 vccd1 _07114_/B sky130_fd_sc_hd__or2_2
XFILLER_0_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_21_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08714_ _08714_/A _08714_/B _08714_/C vssd1 vssd1 vccd1 vccd1 _08717_/B sky130_fd_sc_hd__or3_4
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12914__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ _09692_/B _09692_/C _09692_/A vssd1 vssd1 vccd1 vccd1 _09694_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09791__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ _08546_/X hold2532/X _09222_/B vssd1 vssd1 vccd1 vccd1 _08645_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_156_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout548_A _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13244__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08576_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _08577_/C sky130_fd_sc_hd__xor2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07161__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12287__B _13460_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09999__A1 _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__B _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07527_ hold701/X _13698_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 hold702/A sky130_fd_sc_hd__mux2_1
XFILLER_0_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09999__B2 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__A1 _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ hold278/X _12482_/A vssd1 vssd1 vccd1 vccd1 _14088_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08781__A _08901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13399__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13547__A2 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14933__D _14933_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07389_ _07879_/A _12379_/A _07344_/X vssd1 vssd1 vccd1 vccd1 _07389_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09128_ _09127_/B _09127_/C _09127_/A vssd1 vssd1 vccd1 vccd1 _09129_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_103_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12850__S0 _12950_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ _09056_/A _09057_/Y _08940_/B _08940_/Y vssd1 vssd1 vccd1 vccd1 _09060_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08005__B _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12070_ _14975_/Q _12096_/B _12096_/C _12131_/B vssd1 vssd1 vccd1 vccd1 _12070_/X
+ sky130_fd_sc_hd__or4_1
Xhold570 hold570/A vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 hold581/A vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 hold592/A vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _11201_/B _11019_/X _10797_/X _10802_/B vssd1 vssd1 vccd1 vccd1 _11022_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_109_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _14807_/Q hold683/A _14647_/Q _14743_/Q _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12972_/X sky130_fd_sc_hd__mux4_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1270 _13726_/X vssd1 vssd1 vccd1 vccd1 _15436_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1281 _14302_/Q vssd1 vssd1 vccd1 vccd1 hold1281/X sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ _13744_/A1 hold1105/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11923_/X sky130_fd_sc_hd__mux2_1
X_14711_ _15416_/CLK _14711_/D vssd1 vssd1 vccd1 vccd1 _14711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1292 _07784_/X vssd1 vssd1 vccd1 vccd1 _14399_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _15378_/CLK hold324/X vssd1 vssd1 vccd1 vccd1 hold323/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ hold771/X _13741_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold772/A sky130_fd_sc_hd__mux2_1
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07071__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10805_ _10807_/D vssd1 vssd1 vccd1 vccd1 _10805_/Y sky130_fd_sc_hd__inv_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14573_ _15188_/CLK hold284/X vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_1
X_11785_ hold1505/X _13705_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 _11785_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13524_ _13738_/A1 hold1321/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13524_/X sky130_fd_sc_hd__mux2_1
X_10736_ _10736_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10736_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13455_ _13455_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _15221_/D sky130_fd_sc_hd__and2_1
XFILLER_0_24_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _10666_/B _10666_/C _10666_/A vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11321__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ _07974_/B _08636_/A _13143_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12407_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13102__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ _13386_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _15177_/D sky130_fd_sc_hd__and2_1
X_10598_ _13743_/A1 _11514_/A2 _11514_/B1 _13198_/B _10596_/Y vssd1 vssd1 vccd1 vccd1
+ _10598_/X sky130_fd_sc_hd__a221o_1
X_15125_ _15127_/CLK _15125_/D vssd1 vssd1 vccd1 vccd1 _15125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12337_ hold853/A _13927_/Q _15428_/Q hold2803/X _12466_/S _12343_/A vssd1 vssd1
+ vccd1 vccd1 _12337_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15056_ _15056_/CLK _15056_/D vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__dfxtp_1
X_12268_ _13150_/A _12268_/B vssd1 vssd1 vccd1 vccd1 _14917_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14007_ _15276_/CLK hold292/X vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__dfxtp_1
X_11219_ _11331_/A _11217_/Y _11027_/A _11027_/Y vssd1 vssd1 vccd1 vccd1 _11220_/D
+ sky130_fd_sc_hd__a211o_1
X_12199_ _12211_/S1 _12198_/X _12243_/A vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07925__B1 _11104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11991__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ _14909_/CLK _14909_/D vssd1 vssd1 vccd1 vccd1 hold245/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08585__B _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08350__B1 _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08430_ hold2767/X _08429_/Y _12256_/A vssd1 vssd1 vccd1 vccd1 _08430_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_176_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08361_ _08873_/A _08361_/B vssd1 vssd1 vccd1 vccd1 _08361_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13711__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ _09619_/B _07312_/B vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _08893_/A _09008_/A _08809_/B _08809_/D vssd1 vssd1 vccd1 vccd1 _08294_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07243_ _07241_/Y _07243_/B vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_144_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08405__A1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07174_ _13675_/A1 hold1639/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07174_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08106__A _08107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12851__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout498_A _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12062__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__D _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07156__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08479__C _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 _12953_/B1 vssd1 vssd1 vccd1 vccd1 _13078_/B1 sky130_fd_sc_hd__buf_8
Xfanout368 _07900_/Y vssd1 vssd1 vccd1 vccd1 _12259_/A1 sky130_fd_sc_hd__buf_8
Xfanout379 _12329_/B vssd1 vssd1 vccd1 vccd1 _13103_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09746_ _09745_/A _09745_/B _09745_/C _09745_/D vssd1 vssd1 vccd1 vccd1 _09746_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06958_ _06950_/C _06962_/C _06956_/X _06957_/X vssd1 vssd1 vccd1 vccd1 _06958_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06995__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08776__A _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12899__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09677_ _10185_/A _09979_/C _09678_/C _09824_/A vssd1 vssd1 vccd1 vccd1 _09679_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14928__D _14928_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout832_A _12964_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__B _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__B1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08628_/A vssd1 vssd1 vccd1 vccd1 _08629_/B sky130_fd_sc_hd__inv_2
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ _08989_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _08559_/Y sky130_fd_sc_hd__nor2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _11570_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08644__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _11567_/A _15222_/Q _10522_/A vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__and3_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10451__A1 _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12237__S _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12728__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ _13240_/A _15348_/Q _13240_/C _13241_/D vssd1 vssd1 vccd1 vccd1 fanout6/A
+ sky130_fd_sc_hd__and4_4
XFILLER_0_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _10452_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__or2_1
XFILLER_0_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08016__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12823__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13171_ _13171_/A _13171_/B vssd1 vssd1 vccd1 vccd1 _15036_/D sky130_fd_sc_hd__nor2_1
X_10383_ _10379_/Y _10381_/X _10164_/X _10206_/X vssd1 vssd1 vccd1 vccd1 _10383_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10754__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12122_ _15001_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12122_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13576__B _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12053_ _12059_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _14839_/D sky130_fd_sc_hd__and2_1
XANTENNA__07066__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__xor2_2
Xfanout880 _13360_/A vssd1 vssd1 vccd1 vccd1 _13369_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout891 _13317_/A vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__buf_2
XANTENNA__13000__S0 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__A2 _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08558__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ _12327_/A _12954_/X _12952_/X vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _13661_/A1 hold967/X _11911_/S vssd1 vssd1 vccd1 vccd1 hold968/A sky130_fd_sc_hd__mux2_1
XFILLER_0_158_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12001__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ _12917_/A1 _12885_/X _13050_/S0 vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__a21o_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14625_ _15265_/CLK hold522/X vssd1 vssd1 vccd1 vccd1 hold521/A sky130_fd_sc_hd__dfxtp_1
X_11837_ hold1099/X _13724_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 _11837_/X sky130_fd_sc_hd__mux2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13531__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__S0 _11316_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12967__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14556_ _15421_/CLK _14556_/D vssd1 vssd1 vccd1 vccd1 _14556_/Q sky130_fd_sc_hd__dfxtp_1
X_11768_ hold861/X _13655_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 hold862/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10719_ _10675_/Y _10676_/X _10719_/C _10719_/D vssd1 vssd1 vccd1 vccd1 _10719_/X
+ sky130_fd_sc_hd__and4bb_2
X_13507_ _13721_/A1 hold2011/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13507_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ _15418_/CLK _14487_/D vssd1 vssd1 vccd1 vccd1 _14487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10456__A _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ hold1753/X _13653_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11699_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13438_ _13440_/S _13438_/B vssd1 vssd1 vccd1 vccd1 _13438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12814__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12195__A1 _12128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11986__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10606__D _14966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13369_ _13369_/A _13369_/B vssd1 vssd1 vccd1 vccd1 _15160_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_122_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _15116_/CLK _15108_/D vssd1 vssd1 vccd1 vccd1 _15108_/Q sky130_fd_sc_hd__dfxtp_1
X_07930_ _08201_/A _07929_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_54_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15039_ _15360_/CLK _15039_/D vssd1 vssd1 vccd1 vccd1 hold479/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2707 _10741_/X vssd1 vssd1 vccd1 vccd1 _13400_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2718 _14827_/Q vssd1 vssd1 vccd1 vccd1 hold2718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2729 _15170_/Q vssd1 vssd1 vccd1 vccd1 hold2729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ _15345_/Q _15344_/Q vssd1 vssd1 vccd1 vccd1 _07862_/D sky130_fd_sc_hd__nor2_1
X_09600_ _09599_/B _09599_/C _09599_/A vssd1 vssd1 vccd1 vccd1 _09601_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__11170__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13706__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12610__S _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07792_ hold969/X _13730_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold970/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ _09530_/A _09530_/B _09530_/C vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2797_A _10566_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _09461_/A _09461_/B _09461_/C _09461_/D vssd1 vssd1 vccd1 vccd1 _09464_/C
+ sky130_fd_sc_hd__a22o_1
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08413_ _08413_/A _08474_/A _08413_/C vssd1 vssd1 vccd1 vccd1 _08512_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _09393_/A _09393_/B vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11305__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08344_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08344_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09858__C _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ hold461/A hold733/A hold409/A _14114_/Q _08275_/S0 _07815_/A vssd1 vssd1
+ vccd1 vccd1 _08276_/B sky130_fd_sc_hd__mux4_1
XANTENNA_fanout413_A _06978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__S0 _13066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10984__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ _15202_/Q _11517_/A vssd1 vssd1 vccd1 vccd1 _07227_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11896__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07157_ _13691_/A1 hold1459/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07157_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13396__B _13396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ _13724_/A1 hold2057/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07088_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__C1 _12258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_1__f_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_7_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12894__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07614__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09729_ _09729_/A _09729_/B vssd1 vssd1 vccd1 vccd1 _09731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12740_ hold977/X _14123_/Q _12741_/S vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__mux2_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ hold581/A _15275_/Q _15083_/Q _14376_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12671_/X sky130_fd_sc_hd__mux4_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14410_ _14472_/CLK _14410_/D vssd1 vssd1 vccd1 vccd1 _14410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _11588_/A _11537_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/CLK _15390_/D vssd1 vssd1 vccd1 vccd1 _15390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341_ _15438_/CLK hold632/X vssd1 vssd1 vccd1 vccd1 hold631/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _11553_/A _11553_/B vssd1 vssd1 vccd1 vccd1 _11554_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07825__C1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13049__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10504_ _10295_/Y _10332_/X _10502_/Y _10503_/X vssd1 vssd1 vccd1 vccd1 _10548_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14272_ _15364_/CLK _14272_/D vssd1 vssd1 vccd1 vccd1 _14272_/Q sky130_fd_sc_hd__dfxtp_1
X_11484_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _13372_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_150_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12177__A1 hold2553/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13223_ hold689/X _13669_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold690/A sky130_fd_sc_hd__mux2_1
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10435_ _13742_/A1 _11514_/A2 _12259_/A1 _13197_/B _10433_/Y vssd1 vssd1 vccd1 vccd1
+ _10435_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_150_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07053__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _13389_/A _13154_/B vssd1 vssd1 vccd1 vccd1 _15019_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10366_ _10189_/B _10191_/B _10364_/X _10365_/Y vssd1 vssd1 vccd1 vccd1 _10366_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output165_A _15177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ hold2426/X _12129_/A2 _12104_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ hold469/A _13957_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
X_10297_ _11586_/A _11614_/A _10827_/C vssd1 vssd1 vccd1 vccd1 _10297_/X sky130_fd_sc_hd__and3_1
XANTENNA__11137__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12036_ _12102_/A hold2410/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output332_A _14830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13987_ _15421_/CLK _13987_/D vssd1 vssd1 vccd1 vccd1 _13987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09024__B _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _06943_/A _12933_/X _12937_/X _12988_/C1 vssd1 vssd1 vccd1 vccd1 _12945_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _13100_/S0 _12864_/X _12868_/X _06944_/Y vssd1 vssd1 vccd1 vccd1 _12870_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11570__A _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ _15372_/CLK hold614/X vssd1 vssd1 vccd1 vccd1 hold613/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12404__A2 _12325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08084__A2 _08012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ _15367_/CLK hold654/X vssd1 vssd1 vccd1 vccd1 hold653/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10617__C _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A2 _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ hold415/A _14239_/Q _14399_/Q _14111_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08061_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07011_ _14086_/Q _07875_/B _07643_/C vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__or3_4
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08792__B1 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A2 _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ hold2609/X _08526_/B _08958_/X _08961_/X vssd1 vssd1 vccd1 vccd1 _13388_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_0_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12406__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2504 _15108_/Q vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2515 _14435_/Q vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__buf_1
X_07913_ _06907_/A _08036_/S _08637_/B _07911_/X hold2354/X vssd1 vssd1 vccd1 vccd1
+ _13342_/A sky130_fd_sc_hd__o2111a_1
Xhold2526 _15354_/Q vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__clkbuf_4
X_08893_ _08893_/A _09009_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _08895_/D
+ sky130_fd_sc_hd__nand4_2
Xhold2537 _15346_/Q vssd1 vssd1 vccd1 vccd1 _06907_/A sky130_fd_sc_hd__clkbuf_2
Xhold1803 _14468_/Q vssd1 vssd1 vccd1 vccd1 hold1803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2548 _14975_/Q vssd1 vssd1 vccd1 vccd1 hold2548/X sky130_fd_sc_hd__clkbuf_2
Xhold1814 _13705_/X vssd1 vssd1 vccd1 vccd1 _15411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2559 _12276_/B vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10577__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1825 _14000_/Q vssd1 vssd1 vccd1 vccd1 hold1825/X sky130_fd_sc_hd__dlygate4sd3_1
X_07844_ _15344_/Q _06937_/Y _06938_/Y _15345_/Q vssd1 vssd1 vccd1 vccd1 _07844_/X
+ sky130_fd_sc_hd__o22a_1
Xhold1836 _07624_/X vssd1 vssd1 vccd1 vccd1 _14247_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1847 _13976_/Q vssd1 vssd1 vccd1 vccd1 hold1847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1858 _11986_/X vssd1 vssd1 vccd1 vccd1 _14805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1869 _13892_/Q vssd1 vssd1 vccd1 vccd1 hold1869/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07775_ _13680_/A1 hold1345/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07775_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout363_A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09514_ _09514_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09514_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08847__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11300__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ _10115_/A _09726_/B _09445_/C _09579_/A vssd1 vssd1 vccd1 vccd1 _09579_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout530_A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12576__A _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A _15202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09376_ _09361_/Y _09366_/Y _09375_/X _10246_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _09377_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_164_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08327_ _08420_/A _08327_/B _08327_/C vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__or3_1
XFILLER_0_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10096__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08258_ _08352_/C vssd1 vssd1 vccd1 vccd1 _08258_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12159__A1 hold2538/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ hold2271/X hold2765/A _07214_/S vssd1 vssd1 vccd1 vccd1 _07209_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10824__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__S _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08189_ _08201_/A _08188_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__o21a_1
X_10220_ _10266_/B _10220_/B _10220_/C vssd1 vssd1 vccd1 vccd1 _10220_/X sky130_fd_sc_hd__or3_1
XANTENNA__07609__S _07609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__A1_N _08345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13200__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10151_ _10152_/A _10152_/B _10152_/C vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput280 _14905_/Q vssd1 vssd1 vccd1 vccd1 out0[28] sky130_fd_sc_hd__buf_12
Xoutput291 _14886_/Q vssd1 vssd1 vccd1 vccd1 out0[9] sky130_fd_sc_hd__buf_12
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10082_ _13580_/A _10082_/B vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12331__A1 _13172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ _15443_/CLK _13910_/D vssd1 vssd1 vccd1 vccd1 _13910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14890_ _14987_/CLK _14890_/D vssd1 vssd1 vccd1 vccd1 _14890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__A _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _15080_/CLK hold688/X vssd1 vssd1 vccd1 vccd1 hold687/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12619__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13772_ hold283/X vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__clkbuf_1
X_10984_ _11573_/A _11569_/B _11563_/B _11590_/A vssd1 vssd1 vccd1 vccd1 _10987_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12723_ hold283/A _14314_/Q hold585/A _13974_/Q _12791_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12723_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08683__B _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12654_ _13387_/B _12325_/B _12653_/X vssd1 vssd1 vccd1 vccd1 _12654_/X sky130_fd_sc_hd__a21o_1
X_15442_ _15442_/CLK hold882/X vssd1 vssd1 vccd1 vccd1 hold881/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13044__C1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _11605_/A _11605_/B vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15373_ _15373_/CLK hold846/X vssd1 vssd1 vccd1 vccd1 hold845/A sky130_fd_sc_hd__dfxtp_1
X_12585_ _14664_/Q _13937_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12585_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11536_ _11536_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__nand2_1
X_14324_ _15416_/CLK hold962/X vssd1 vssd1 vccd1 vccd1 hold961/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output282_A _14879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14255_ _15090_/CLK _14255_/D vssd1 vssd1 vccd1 vccd1 _14255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11467_ _11467_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07519__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ hold2227/X _13652_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13206_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09566__A2 _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10418_ _15383_/Q _15286_/Q hold393/A _14387_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10418_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09110__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14186_ _15278_/CLK hold178/X vssd1 vssd1 vccd1 vccd1 _14186_/Q sky130_fd_sc_hd__dfxtp_1
X_11398_ _11626_/B _11397_/B _11397_/C vssd1 vssd1 vccd1 vccd1 _11399_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13137_ _13495_/A hold141/X vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__and2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10350_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10349_/Y sky130_fd_sc_hd__nor2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A1 _13065_/X _13067_/X vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12322__A1 _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _12059_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _14822_/D sky130_fd_sc_hd__and2_1
XFILLER_0_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11530__C1 _15227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07560_ _13393_/A hold125/X vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__and2_1
XFILLER_0_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07491_ hold1727/X _13730_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07491_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ _09941_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09161_ _09162_/A _09162_/B vssd1 vssd1 vccd1 vccd1 _09161_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08112_ _08050_/X _08111_/X _08441_/B vssd1 vssd1 vccd1 vccd1 _08112_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11061__A1 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09092_ _11104_/A _12275_/B _09091_/X vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08043_ _08049_/B vssd1 vssd1 vccd1 vccd1 _08043_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold900 hold900/A vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold911 hold911/A vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold922 hold922/A vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A0 hold2621/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__S0 _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold933 hold933/A vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 hold944/A vssd1 vssd1 vccd1 vccd1 hold944/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08114__A _14430_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold955 hold955/A vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 hold966/A vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 hold977/A vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _09993_/B _09993_/C _09993_/A vssd1 vssd1 vccd1 vccd1 _09995_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold988 hold988/A vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 hold999/A vssd1 vssd1 vccd1 vccd1 hold999/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07953__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2301 _14482_/Q vssd1 vssd1 vccd1 vccd1 hold2301/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2312 _14056_/Q vssd1 vssd1 vccd1 vccd1 _07852_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08945_ _08944_/B _08944_/C _08944_/A vssd1 vssd1 vccd1 vccd1 _08945_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2323 _12181_/X vssd1 vssd1 vccd1 vccd1 _14901_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout480_A _06959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2334 _13425_/X vssd1 vssd1 vccd1 vccd1 _15206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1600 _07539_/X vssd1 vssd1 vccd1 vccd1 _14164_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2345 _14031_/Q vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout578_A _07448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2356 _13750_/B vssd1 vssd1 vccd1 vccd1 _13341_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1611 _15281_/Q vssd1 vssd1 vccd1 vccd1 hold1611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2367 _13752_/X vssd1 vssd1 vccd1 vccd1 _15459_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08876_ hold791/A _13940_/Q _15441_/Q _13908_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _08877_/B sky130_fd_sc_hd__mux4_1
Xhold1622 _07604_/X vssd1 vssd1 vccd1 vccd1 _14228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1633 _14544_/Q vssd1 vssd1 vccd1 vccd1 hold1633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2378 _07969_/Y vssd1 vssd1 vccd1 vccd1 _13412_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2389 _13597_/X vssd1 vssd1 vccd1 vccd1 _15324_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 _13688_/X vssd1 vssd1 vccd1 vccd1 _15394_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07164__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1655 _15434_/Q vssd1 vssd1 vccd1 vccd1 hold1655/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__B _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ hold525/A hold327/A _14396_/Q hold517/A _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _07828_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1666 _07589_/X vssd1 vssd1 vccd1 vccd1 _14213_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1677 _13950_/Q vssd1 vssd1 vccd1 vccd1 hold1677/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07740__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1688 _07040_/X vssd1 vssd1 vccd1 vccd1 _13857_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1699 _13915_/Q vssd1 vssd1 vccd1 vccd1 hold1699/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07758_ _13663_/A1 hold1829/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07758_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14936__D _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ hold817/X _13662_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold818/A sky130_fd_sc_hd__mux2_1
XANTENNA__09493__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _10129_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ _13880_/Q _14008_/Q hold663/A _13816_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09359_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_165_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12475__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12370_ _12692_/A1 _12369_/X _12368_/X _12669_/A1 vssd1 vssd1 vccd1 vccd1 _12370_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08453__C1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ hold2786/X input24/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_132_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07008__A0 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _14042_/CLK _14040_/D vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ _11252_/A _11252_/B _11252_/C vssd1 vssd1 vccd1 vccd1 _11254_/B sky130_fd_sc_hd__nand3_2
XANTENNA__08205__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10238__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ _09993_/B _09995_/B _10201_/X _10202_/Y vssd1 vssd1 vccd1 vccd1 _10206_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09953__C1 _11511_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _11183_/A _11183_/B _11371_/B _11183_/D vssd1 vssd1 vccd1 vccd1 _11183_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _10306_/A _11168_/A _10135_/C _10135_/D vssd1 vssd1 vccd1 vccd1 _10134_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_101_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13584__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10065_ _10065_/A _10065_/B _10065_/C vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__nand3_1
X_14942_ _15293_/CLK _14942_/D vssd1 vssd1 vccd1 vccd1 _14942_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__10315__B1 _14957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ _14876_/CLK _14873_/D vssd1 vssd1 vccd1 vccd1 _14873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15007__D _15007_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13824_ _14791_/CLK _13824_/D vssd1 vssd1 vccd1 vccd1 _13824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07802__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10618__A1 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10967_ _11596_/A _11597_/A _11573_/B _14966_/Q vssd1 vssd1 vccd1 vccd1 _11150_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08287__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13755_ hold2632/X _07926_/A _13754_/X _13409_/A vssd1 vssd1 vccd1 vccd1 _13755_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_202_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _13106_/A1 _13155_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12707_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10898_ _10713_/B _10713_/Y _10896_/A _10897_/X vssd1 vssd1 vccd1 vccd1 _11089_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13686_ hold1163/X hold479/X _13698_/S vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10448__B _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15425_ _15425_/CLK _15425_/D vssd1 vssd1 vccd1 vccd1 _15425_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_31_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12637_ _12689_/S1 _12634_/X _12636_/X vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11043__A1 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15356_ _15356_/CLK _15356_/D vssd1 vssd1 vccd1 vccd1 _15356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12568_ _12368_/A _12565_/X _12567_/X vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06942__A _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11519_ _11383_/A _11383_/B _11384_/Y vssd1 vssd1 vccd1 vccd1 _11521_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14307_ _15270_/CLK _14307_/D vssd1 vssd1 vccd1 vccd1 _14307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ _13869_/Q hold717/A _13837_/Q hold745/A _12460_/S _12689_/S1 vssd1 vssd1
+ vccd1 vccd1 _12499_/X sky130_fd_sc_hd__mux4_1
X_15287_ _15287_/CLK hold450/X vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__dfxtp_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _15434_/CLK _14238_/D vssd1 vssd1 vccd1 vccd1 _14238_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09095__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10183__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08747__B1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__A1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09972__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ _15418_/CLK _14169_/D vssd1 vssd1 vccd1 vccd1 _14169_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08211__A2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08869__A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 _15042_/Q vssd1 vssd1 vccd1 vccd1 _13689_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _13663_/A1 hold1305/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06991_/X sky130_fd_sc_hd__mux2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2410_A _14831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08727_/Y _08728_/X _08621_/Y _08623_/Y vssd1 vssd1 vccd1 vccd1 _08731_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ hold997/A _13938_/Q hold955/A _13906_/Q _08763_/S0 _08763_/S1 vssd1 vssd1
+ vccd1 vccd1 _08662_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07612_ hold2085/X _13718_/A1 _07626_/S vssd1 vssd1 vccd1 vccd1 _07612_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13714__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08592_ _08592_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07712__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07543_ hold357/X _13714_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold358/A sky130_fd_sc_hd__mux2_1
XANTENNA__10639__A _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07474_ hold267/X _07474_/B vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__and2_1
XFILLER_0_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10358__B _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09213_ _09214_/B _09213_/B vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09227__A1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09144_ _09145_/A _09145_/B vssd1 vssd1 vccd1 vccd1 _09146_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_161_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ _09075_/A _09075_/B _09075_/C vssd1 vssd1 vccd1 vccd1 _09075_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12209__S1 _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08026_ _12256_/A _12258_/S vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__nand2_8
XANTENNA__07159__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1 fanout2/A vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__buf_4
XANTENNA__11189__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold730 hold730/A vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 hold741/A vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 hold752/A vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 hold763/A vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06998__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 hold774/A vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 hold785/A vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 hold796/A vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09977_ _09860_/A _09860_/B _09857_/X _09858_/X _09709_/B vssd1 vssd1 vccd1 vccd1
+ _09982_/A sky130_fd_sc_hd__a32o_1
XANTENNA_fanout862_A _06946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2120 _07764_/X vssd1 vssd1 vccd1 vccd1 _14380_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2131 _15366_/Q vssd1 vssd1 vccd1 vccd1 hold2131/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2142 _07747_/X vssd1 vssd1 vccd1 vccd1 _14363_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _08928_/A _09039_/B _08928_/C vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__nand3_2
Xhold2153 _13885_/Q vssd1 vssd1 vccd1 vccd1 hold2153/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2164 _11734_/X vssd1 vssd1 vccd1 vccd1 _14528_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2175 _13865_/Q vssd1 vssd1 vccd1 vccd1 hold2175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 _07675_/X vssd1 vssd1 vccd1 vccd1 _14296_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2186 _07103_/X vssd1 vssd1 vccd1 vccd1 _13916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _14264_/Q vssd1 vssd1 vccd1 vccd1 hold1441/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2197 _14718_/Q vssd1 vssd1 vccd1 vccd1 hold2197/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _07212_/X vssd1 vssd1 vccd1 vccd1 _14019_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1463 _14361_/Q vssd1 vssd1 vccd1 vccd1 hold1463/X sky130_fd_sc_hd__dlygate4sd3_1
X_08859_ _08256_/A _13355_/B _08857_/X _08858_/Y vssd1 vssd1 vccd1 vccd1 _08859_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1474 _13210_/X vssd1 vssd1 vccd1 vccd1 _15074_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 _14206_/Q vssd1 vssd1 vccd1 vccd1 hold1485/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _07000_/X vssd1 vssd1 vccd1 vccd1 _13819_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ hold543/X _13691_/A1 _11877_/S vssd1 vssd1 vccd1 vccd1 hold544/A sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07622__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ _11614_/A _11378_/C _11378_/D _11586_/A vssd1 vssd1 vccd1 vccd1 _10821_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12696__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ _14426_/Q _07919_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13540_/X sky130_fd_sc_hd__mux2_1
X_10752_ _11113_/C vssd1 vssd1 vccd1 vccd1 _10752_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13471_ _13479_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13471_/X sky130_fd_sc_hd__and2_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10683_ _10510_/B _10510_/C _10510_/A vssd1 vssd1 vccd1 vccd1 _10684_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12448__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15210_ _15226_/CLK _15210_/D vssd1 vssd1 vccd1 vccd1 _15210_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12422_ _14785_/Q hold483/A hold521/A _14721_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12422_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_152_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08977__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12353_ _12352_/X hold2804/X _12601_/A vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__mux2_1
X_15141_ _15304_/CLK _15141_/D vssd1 vssd1 vccd1 vccd1 _15141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07069__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11304_ _11507_/A _11301_/X _11303_/X vssd1 vssd1 vccd1 vccd1 _11304_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15072_ _15072_/CLK hold936/X vssd1 vssd1 vccd1 vccd1 hold935/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12284_ _13479_/A _12284_/B vssd1 vssd1 vccd1 vccd1 _14933_/D sky130_fd_sc_hd__and2_2
XFILLER_0_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ _15293_/CLK _14023_/D vssd1 vssd1 vccd1 vccd1 _14023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11235_ _11047_/B _11049_/B _11047_/A vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11166_ _11569_/A _11605_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11166_/X sky130_fd_sc_hd__and3_1
XFILLER_0_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07952__A1 _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10117_ _10115_/X _10117_/B vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07952__B2 _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _11098_/A _11098_/B _11096_/Y vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_93_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12828__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10839__A1 _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ _09885_/Y _09887_/X _10046_/X _10047_/Y vssd1 vssd1 vccd1 vccd1 _10050_/B
+ sky130_fd_sc_hd__o211ai_4
X_14925_ _15247_/CLK _14925_/D vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10839__B2 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08052__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13534__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10934__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14856_ _15004_/CLK _14856_/D vssd1 vssd1 vccd1 vccd1 _14856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07532__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13807_ _15391_/CLK _13807_/D vssd1 vssd1 vccd1 vccd1 _13807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10459__A _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14787_ _15299_/CLK _14787_/D vssd1 vssd1 vccd1 vccd1 _14787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _14095_/Q _12131_/A _14097_/Q _14096_/Q vssd1 vssd1 vccd1 vccd1 _12056_/S
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13738_ hold1119/X _13738_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12461__B1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__B _15220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__S _11993_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09967__B _10338_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13669_ hold1867/X _13669_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 _13669_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12439__S1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _15408_/CLK _15408_/D vssd1 vssd1 vccd1 vccd1 _15408_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11016__B2 _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ hold717/X _13691_/A1 _07198_/S vssd1 vssd1 vccd1 vccd1 hold718/A sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ _15357_/CLK _15339_/D vssd1 vssd1 vccd1 vccd1 _15339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08432__A2 _13383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _09693_/Y _09696_/Y _09898_/Y _09899_/X vssd1 vssd1 vccd1 vccd1 _09900_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__13709__S _13714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B1 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout506 _06926_/Y vssd1 vssd1 vccd1 vccd1 _12201_/C1 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07707__S _07709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ _09831_/A _09831_/B _09831_/C vssd1 vssd1 vccd1 vccd1 _09833_/B sky130_fd_sc_hd__nand3_2
Xfanout517 _12241_/A vssd1 vssd1 vccd1 vccd1 _08760_/A sky130_fd_sc_hd__clkbuf_8
Xfanout528 _15425_/Q vssd1 vssd1 vccd1 vccd1 _10255_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout539 _08763_/S1 vssd1 vssd1 vccd1 vccd1 _08130_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_193_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ _09762_/A _09762_/B _09762_/C _09759_/X vssd1 vssd1 vccd1 vccd1 _09763_/B
+ sky130_fd_sc_hd__or4b_2
X_06974_ _14093_/Q _14092_/Q _06973_/X _06972_/X vssd1 vssd1 vccd1 vccd1 _07643_/C
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08713_ _08712_/B _08712_/C _08712_/A vssd1 vssd1 vccd1 vccd1 _08714_/C sky130_fd_sc_hd__a21oi_1
X_09693_ _09693_/A vssd1 vssd1 vccd1 vccd1 _09693_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08644_ _09918_/A _13428_/B _08643_/X _10233_/A vssd1 vssd1 vccd1 vccd1 _08644_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09791__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08575_ _09858_/A _08574_/X _08573_/X vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__a21bo_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout443_A _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ hold1065/X _13730_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07526_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11899__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ _07457_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14087_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout610_A _15207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08781__B _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07388_ _07879_/A _12379_/A _07344_/X vssd1 vssd1 vccd1 vccd1 _07981_/A sky130_fd_sc_hd__o21a_2
XANTENNA__13399__B _13399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ _09127_/A _09127_/B _09127_/C vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__nor3_1
XANTENNA__12755__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12850__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09058_ _08940_/B _08940_/Y _09056_/A _09057_/Y vssd1 vssd1 vccd1 vccd1 _09060_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08009_ _08010_/A _08010_/B _08010_/C vssd1 vssd1 vccd1 vccd1 _08009_/X sky130_fd_sc_hd__and3_1
XANTENNA__08005__C _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold560 hold560/A vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 hold571/A vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _10797_/X _10802_/B _11201_/B _11019_/X vssd1 vssd1 vccd1 vccd1 _11022_/B
+ sky130_fd_sc_hd__o211ai_2
Xhold582 hold582/A vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07617__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold593 hold593/A vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11139__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ hold315/A hold449/X hold523/A hold1781/X _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12971_/X sky130_fd_sc_hd__mux4_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1260 _13220_/X vssd1 vssd1 vccd1 vccd1 _15084_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1271 _14487_/Q vssd1 vssd1 vccd1 vccd1 hold1271/X sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ _15452_/CLK hold332/X vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__dfxtp_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1282 _07682_/X vssd1 vssd1 vccd1 vccd1 _14302_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ hold2765/A hold1903/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__mux2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1293 _14225_/Q vssd1 vssd1 vccd1 vccd1 hold1293/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _15376_/CLK hold616/X vssd1 vssd1 vccd1 vccd1 hold615/A sky130_fd_sc_hd__dfxtp_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ hold607/X _13740_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold608/A sky130_fd_sc_hd__mux2_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11246__A1 _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _11598_/A _11590_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _10807_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_83_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _15179_/CLK hold250/X vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dfxtp_1
X_11784_ hold1909/X _13671_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08111__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08111__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__A1 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13671_/A1 hold1611/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13523_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10735_ _10562_/A _10559_/X _10561_/B vssd1 vssd1 vccd1 vccd1 _10735_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ _10666_/A _10666_/B _10666_/C vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__and3_2
X_13454_ _10405_/B _12284_/B _13468_/A vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output195_A _06963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _12327_/A _12404_/X _12402_/X vssd1 vssd1 vccd1 vccd1 _13143_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_207_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13385_ _13386_/A _13385_/B vssd1 vssd1 vccd1 vccd1 _15176_/D sky130_fd_sc_hd__and2_1
XFILLER_0_140_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10597_ hold2760/X input19/X _12253_/S vssd1 vssd1 vccd1 vccd1 _13198_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15124_ _15132_/CLK _15124_/D vssd1 vssd1 vccd1 vccd1 _15124_/Q sky130_fd_sc_hd__dfxtp_1
X_12336_ hold509/A hold497/X _14139_/Q _14457_/Q _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12336_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_120_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13529__S _13534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055_ _15087_/CLK _15055_/D vssd1 vssd1 vccd1 vccd1 _15055_/Q sky130_fd_sc_hd__dfxtp_1
X_12267_ _13150_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _14916_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ _11027_/A _11027_/Y _11331_/A _11217_/Y vssd1 vssd1 vccd1 vccd1 _11331_/B
+ sky130_fd_sc_hd__o211ai_2
X_14006_ _14472_/CLK _14006_/D vssd1 vssd1 vccd1 vccd1 _14006_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07527__S _07528_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08212__A _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12198_ _14589_/Q _13958_/Q _12198_/S vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07925__B2 _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ _11578_/C _11149_/B vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__A _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _14992_/CLK _14908_/D vssd1 vssd1 vccd1 vccd1 _14908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08585__C _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09043__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14839_ _14842_/CLK _14839_/D vssd1 vssd1 vccd1 vccd1 _14839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ hold665/A _14502_/Q hold569/A _14726_/Q _08868_/S0 _08868_/S1 vssd1 vssd1
+ vccd1 vccd1 _08361_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08882__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ _11378_/D _10283_/C vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__or2_1
X_08291_ _08893_/A _09008_/A _09542_/A _08809_/D vssd1 vssd1 vccd1 vccd1 _08401_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_184_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07242_ _10356_/C _11588_/B vssd1 vssd1 vccd1 vccd1 _07243_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12737__A1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07173_ _13674_/A1 hold1855/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12596__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A _07745_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__C1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09814_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09814_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08479__D _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 _12330_/X vssd1 vssd1 vccd1 vccd1 _12953_/B1 sky130_fd_sc_hd__clkbuf_16
Xfanout369 _12260_/A2 vssd1 vssd1 vccd1 vccd1 _11514_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_94_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09745_ _09745_/A _09745_/B _09745_/C _09745_/D vssd1 vssd1 vccd1 vccd1 _09745_/X
+ sky130_fd_sc_hd__or4_2
X_06957_ _14030_/Q _14036_/Q hold237/A hold273/A vssd1 vssd1 vccd1 vccd1 _06957_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout560_A _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13465__A2 _13468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12899__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _10183_/A _09979_/B _09860_/B _09676_/D vssd1 vssd1 vccd1 vccd1 _09824_/A
+ sky130_fd_sc_hd__nand4_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07172__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__C _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08627_ _08515_/X _08517_/X _08624_/X _08625_/Y vssd1 vssd1 vccd1 vccd1 _08628_/A
+ sky130_fd_sc_hd__o211a_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout825_A _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09888__A _09888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08558_ hold993/A _14213_/Q _14149_/Q _14467_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08559_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13622__C1 _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ hold1921/X _13748_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07509_/X sky130_fd_sc_hd__mux2_1
X_08489_ _09164_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _08491_/C sky130_fd_sc_hd__and2_1
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10827__A _14953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08644__A2 _13428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ _11567_/A _15222_/Q vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13203__A _13404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10451__A2 _11605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10451_ _11598_/A _11605_/B _10450_/C _10450_/D vssd1 vssd1 vccd1 vccd1 _10452_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_162_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08016__B _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12823__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13170_ _13171_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _15035_/D sky130_fd_sc_hd__nor2_1
X_10382_ _10164_/X _10206_/X _10379_/Y _10381_/X vssd1 vssd1 vccd1 vccd1 _10382_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12121_ hold2491/X _12129_/A2 _12120_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12253__S _12253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12052_ hold2535/X hold2716/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12052_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold390 hold390/A vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _11620_/A _11564_/B vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12339__S0 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 _13487_/A vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout881 _13373_/A vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13592__B _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout892 _13317_/A vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__buf_6
XFILLER_0_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13000__S1 _13100_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _10566_/Y _12325_/B _12953_/X vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__a21o_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07082__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 _07023_/X vssd1 vssd1 vccd1 vccd1 _13840_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _13512_/A0 hold1585/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_197_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12885_ hold607/A _13949_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12885_/X sky130_fd_sc_hd__mux2_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _15264_/CLK hold924/X vssd1 vssd1 vccd1 vccd1 hold923/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09798__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11836_ hold2815/X hold465/X _11845_/S vssd1 vssd1 vccd1 vccd1 hold466/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07810__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_97_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__S1 _11316_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12967__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _15287_/CLK _14555_/D vssd1 vssd1 vccd1 vccd1 _14555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11767_ hold971/X _13654_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 hold972/A sky130_fd_sc_hd__mux2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08191__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ _13654_/A1 hold2261/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_140_clk_A clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ _10717_/B _10717_/C _10717_/A vssd1 vssd1 vccd1 vccd1 _10719_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_99_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _14958_/CLK _14486_/D vssd1 vssd1 vccd1 vccd1 _14486_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10456__B _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11698_ hold2067/X _13652_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 _11698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12719__A1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_20_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ _13455_/A _13437_/B vssd1 vssd1 vccd1 vccd1 _15212_/D sky130_fd_sc_hd__and2_1
XFILLER_0_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ _10646_/Y _10647_/X _10473_/X _10476_/X vssd1 vssd1 vccd1 vccd1 _10650_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12952__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__A1 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12814__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13368_ _13369_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _15159_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_155_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ _15116_/CLK _15107_/D vssd1 vssd1 vccd1 vccd1 _15107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12319_ hold165/A hold529/A _14589_/Q _13958_/Q _12466_/S _12365_/S1 vssd1 vssd1
+ vccd1 vccd1 _12319_/X sky130_fd_sc_hd__mux4_1
X_13299_ _13317_/A _13299_/B vssd1 vssd1 vccd1 vccd1 _15119_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_35_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ _15427_/CLK _15038_/D vssd1 vssd1 vccd1 vccd1 _15038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2708 _14815_/Q vssd1 vssd1 vccd1 vccd1 hold2708/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2719 _12028_/X vssd1 vssd1 vccd1 vccd1 _12029_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07860_ _14061_/Q _07343_/X _07859_/Y _07342_/X vssd1 vssd1 vccd1 vccd1 _12379_/B
+ sky130_fd_sc_hd__o211a_2
XANTENNA__08877__A _08877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07791_ hold1865/X _13729_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 _07791_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08596__B _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ _09530_/A _09530_/B _09530_/C vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__and3_1
XFILLER_0_79_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ _09461_/A _09461_/B _09461_/C _09461_/D vssd1 vssd1 vccd1 vccd1 _09464_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__12750__S0 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2692_A _14434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_184_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15040_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13722__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _08411_/A _08468_/B _08411_/C vssd1 vssd1 vccd1 vccd1 _08413_/C sky130_fd_sc_hd__a21o_1
X_09392_ _09392_/A _09392_/B vssd1 vssd1 vccd1 vccd1 _09393_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07720__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ _08255_/A _08252_/Y _08254_/B vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11305__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_clk_A clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07834__B1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _12241_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07225_ _09138_/A _11517_/A vssd1 vssd1 vccd1 vccd1 _08496_/A sky130_fd_sc_hd__and2_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout406_A _07182_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ _13657_/A1 hold2291/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07087_ _13690_/A1 hold2147/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07087_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07167__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07996__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14939__D _14939_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ _08197_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _07989_/X sky130_fd_sc_hd__or2_1
X_09728_ _09729_/B _09729_/A vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12102__A _12102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _10166_/A _10338_/B _09979_/D _09809_/C vssd1 vssd1 vccd1 vccd1 _09813_/A
+ sky130_fd_sc_hd__nand4_2
Xclkbuf_leaf_175_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15268_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_195_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ _12670_/A _12670_/B _12601_/A vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_195_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07630__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__xor2_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08672__D _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14340_ _14956_/CLK hold320/X vssd1 vssd1 vccd1 vccd1 hold319/A sky130_fd_sc_hd__dfxtp_1
X_11552_ _11552_/A _11552_/B vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_108_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13049__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _10502_/A _10502_/B _10502_/C _10502_/D vssd1 vssd1 vccd1 vccd1 _10503_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11483_ _11482_/A _11482_/B _11484_/A vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__a21o_1
X_14271_ _15395_/CLK hold504/X vssd1 vssd1 vccd1 vccd1 hold503/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13222_ hold347/X _13668_/A1 _13236_/S vssd1 vssd1 vccd1 vccd1 hold348/A sky130_fd_sc_hd__mux2_1
X_10434_ hold2695/X input18/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10365_ _10364_/B _10364_/C _10364_/A vssd1 vssd1 vccd1 vccd1 _10365_/Y sky130_fd_sc_hd__a21oi_2
X_13153_ _13389_/A _13153_/B vssd1 vssd1 vccd1 vccd1 _15018_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07077__S _07077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12104_ _14992_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12104_/X
+ sky130_fd_sc_hd__or4_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ hold361/X hold2003/X _13091_/S vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10296_ _10296_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__xor2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12035_ _12037_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _14830_/D sky130_fd_sc_hd__and2_1
XFILLER_0_109_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13108__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ _14483_/CLK _13986_/D vssd1 vssd1 vccd1 vccd1 _13986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12101__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09502__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _13024_/S1 _12934_/X _12936_/X vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_166_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _14409_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12868_ _13074_/S1 _12865_/X _12867_/X vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07540__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__B _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607_ _15374_/CLK hold542/X vssd1 vssd1 vccd1 vccd1 hold541/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ hold2065/X _13673_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13601__A2 _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ _13881_/Q _14009_/Q hold565/A _13817_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12799_/X sky130_fd_sc_hd__mux4_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14538_ _15438_/CLK _14538_/D vssd1 vssd1 vccd1 vccd1 _14538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10617__D _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12682__A _13150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469_ _14602_/CLK _14469_/D vssd1 vssd1 vccd1 vccd1 _14469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07010_ _13748_/A1 hold1409/X _07010_/S vssd1 vssd1 vccd1 vccd1 _07010_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12799__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2538_A _14986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08792__A1 _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08792__B2 _08908_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _08960_/X _09075_/C vssd1 vssd1 vccd1 vccd1 _08961_/X sky130_fd_sc_hd__and2b_1
Xhold2505 _08250_/B vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13717__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07912_ _06907_/A _08036_/S _07911_/X vssd1 vssd1 vccd1 vccd1 _07912_/X sky130_fd_sc_hd__o21a_1
Xhold2516 _15171_/Q vssd1 vssd1 vccd1 vccd1 hold2516/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2527 _15164_/Q vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08892_ _08892_/A _09008_/A _09864_/C _09864_/D vssd1 vssd1 vccd1 vccd1 _08892_/X
+ sky130_fd_sc_hd__and4_1
Xhold2538 _14986_/Q vssd1 vssd1 vccd1 vccd1 hold2538/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1804 _11665_/X vssd1 vssd1 vccd1 vccd1 _14468_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07715__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2549 _12137_/X vssd1 vssd1 vccd1 vccd1 _14879_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1815 _13946_/Q vssd1 vssd1 vccd1 vccd1 hold1815/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12971__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ _15342_/Q _06935_/Y _07838_/Y _07842_/X _15293_/Q vssd1 vssd1 vccd1 vccd1
+ _07843_/X sky130_fd_sc_hd__o2111a_1
Xhold1826 _07193_/X vssd1 vssd1 vccd1 vccd1 _14000_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08400__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1837 _14292_/Q vssd1 vssd1 vccd1 vccd1 hold1837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1848 _07168_/X vssd1 vssd1 vccd1 vccd1 _13976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1859 _13876_/Q vssd1 vssd1 vccd1 vccd1 hold1859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _13679_/A1 hold1535/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07774_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12723__S0 _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ hold721/A _13945_/Q hold511/A _13913_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09514_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_157_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _15395_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10103__A1 _11510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ _10002_/C _10110_/A _09724_/C _09724_/D vssd1 vssd1 vccd1 vccd1 _09579_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ _10255_/A1 _09368_/Y _09370_/Y _09372_/Y _09374_/Y vssd1 vssd1 vccd1 vccd1
+ _09375_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13053__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout523_A _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08326_ _08162_/A _08326_/B vssd1 vssd1 vccd1 vccd1 _08327_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ _08257_/A _14430_/Q _08257_/C vssd1 vssd1 vccd1 vccd1 _08352_/C sky130_fd_sc_hd__and3_1
XFILLER_0_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11700__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ hold1503/X _13742_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 _07208_/X sky130_fd_sc_hd__mux2_1
X_08188_ _13869_/Q hold717/A _13837_/Q hold745/A _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08188_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout892_A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__B _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07139_ _13740_/A1 hold1965/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13200__B _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11001__A _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10150_ _10038_/A _10038_/C _10038_/B vssd1 vssd1 vccd1 vccd1 _10152_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput270 _14896_/Q vssd1 vssd1 vccd1 vccd1 out0[19] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput281 _14906_/Q vssd1 vssd1 vccd1 vccd1 out0[29] sky130_fd_sc_hd__buf_12
Xoutput292 _14845_/Q vssd1 vssd1 vccd1 vccd1 out1[0] sky130_fd_sc_hd__buf_12
X_10081_ _13749_/A _13450_/B vssd1 vssd1 vccd1 vccd1 _10081_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12867__B1 _14490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__S _07626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__A2 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09125__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _15079_/CLK _13840_/D vssd1 vssd1 vccd1 vccd1 _13840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12714__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ hold249/X vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_148_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15416_/CLK sky130_fd_sc_hd__clkbuf_16
X_10983_ _10983_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ _14797_/Q _14509_/Q _14637_/Q _14733_/Q _12741_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12722_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_167_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11390__B _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15441_ _15441_/CLK _15441_/D vssd1 vssd1 vccd1 vccd1 _15441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _13664_/A1 _12329_/B _12953_/B1 _13185_/B vssd1 vssd1 vccd1 vccd1 _12653_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11604_ _11604_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ _15372_/CLK hold582/X vssd1 vssd1 vccd1 vccd1 hold581/A sky130_fd_sc_hd__dfxtp_1
X_12584_ _15438_/Q _13905_/Q _12591_/S vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14323_ _15382_/CLK hold628/X vssd1 vssd1 vccd1 vccd1 hold627/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11535_ _11535_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14254_ _15089_/CLK hold534/X vssd1 vssd1 vccd1 vccd1 hold533/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _11466_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11467_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09646__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ hold1039/X _13651_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10417_ _15424_/Q _10414_/X _10416_/X vssd1 vssd1 vccd1 vccd1 _10417_/Y sky130_fd_sc_hd__o21ai_1
X_11397_ _11626_/B _11397_/B _11397_/C vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__nand3_1
X_14185_ _15184_/CLK hold126/X vssd1 vssd1 vccd1 vccd1 _14185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12007__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _13499_/A hold101/X vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__and2_1
X_10348_ _10175_/A _10174_/Y _10171_/X vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__xnor2_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12441__S _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ _13092_/A1 _13066_/X _06943_/A vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10750__A _13750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09723__B1 _09724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ hold2607/X hold2686/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12019_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08220__A _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11530__B1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13969_ _15268_/CLK _13969_/D vssd1 vssd1 vccd1 vccd1 _13969_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_139_clk clkbuf_4_9__f_clk/X vssd1 vssd1 vccd1 vccd1 _15380_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12677__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07490_ hold1527/X _13729_/A1 _07493_/S vssd1 vssd1 vccd1 vccd1 _07490_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_159_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09703__A1_N _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ _09160_/A _09160_/B vssd1 vssd1 vccd1 vccd1 _09162_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08111_ _09918_/A _13416_/B _13347_/B _08256_/A _08110_/Y vssd1 vssd1 vccd1 vccd1
+ _08111_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_173_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12794__C1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09091_ _08256_/A _13357_/B _09089_/X _09090_/Y vssd1 vssd1 vccd1 vccd1 _09091_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11061__A2 _11620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12616__S _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__B1 _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _14428_/Q _08042_/B _14426_/Q vssd1 vssd1 vccd1 vccd1 _08049_/B sky130_fd_sc_hd__and3_1
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09637__S0 _09795_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 hold901/A vssd1 vssd1 vccd1 vccd1 hold901/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold912 hold912/A vssd1 vssd1 vccd1 vccd1 hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 hold923/A vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 hold934/A vssd1 vssd1 vccd1 vccd1 hold934/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10247__S1 _10425_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 hold945/A vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 hold956/A vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 hold967/A vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 hold978/A vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _09993_/A _09993_/B _09993_/C vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_12_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold989 hold989/A vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2302 _11679_/X vssd1 vssd1 vccd1 vccd1 _14482_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ _08944_/A _08944_/B _08944_/C vssd1 vssd1 vccd1 vccd1 _08944_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__07953__B _08892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2313 _14026_/Q vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2324 hold2827/X vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__buf_1
XFILLER_0_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2335 _14913_/Q vssd1 vssd1 vccd1 vccd1 _13474_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2346 _15309_/Q vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__buf_1
Xhold1601 _15386_/Q vssd1 vssd1 vccd1 vccd1 hold1601/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1612 _13523_/X vssd1 vssd1 vccd1 vccd1 _15281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2357 _15160_/Q vssd1 vssd1 vccd1 vccd1 hold2357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1623 _14472_/Q vssd1 vssd1 vccd1 vccd1 hold1623/X sky130_fd_sc_hd__dlygate4sd3_1
X_08875_ _08877_/A _08875_/B vssd1 vssd1 vccd1 vccd1 _08875_/Y sky130_fd_sc_hd__nor2_1
Xhold2368 _15331_/Q vssd1 vssd1 vccd1 vccd1 _06913_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1634 _11750_/X vssd1 vssd1 vccd1 vccd1 _14544_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2379 hold2849/X vssd1 vssd1 vccd1 vccd1 _08535_/B sky130_fd_sc_hd__buf_1
XFILLER_0_93_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1645 _14149_/Q vssd1 vssd1 vccd1 vccd1 hold1645/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1656 _13724_/X vssd1 vssd1 vccd1 vccd1 _15434_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07826_ _12241_/A _07826_/B vssd1 vssd1 vccd1 vccd1 _07826_/Y sky130_fd_sc_hd__nor2_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__C _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1667 _13912_/Q vssd1 vssd1 vccd1 vccd1 hold1667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1678 _07140_/X vssd1 vssd1 vccd1 vccd1 _13950_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1689 _13803_/Q vssd1 vssd1 vccd1 vccd1 hold1689/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout640_A _15200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ _13662_/A1 hold1709/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07757_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10088__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11824__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07688_ hold505/X _13661_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold506/A sky130_fd_sc_hd__mux2_1
XANTENNA__09493__A2 _13442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09427_ _10010_/B _09427_/B vssd1 vssd1 vccd1 vccd1 _09587_/A sky130_fd_sc_hd__and2_2
XFILLER_0_137_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08128__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09358_ hold239/A _14316_/Q hold541/A _13976_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09358_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09245__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08309_ _08310_/A _08310_/B _08310_/C vssd1 vssd1 vccd1 vccd1 _08309_/X sky130_fd_sc_hd__and3_1
XFILLER_0_180_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09289_ _09288_/A _09288_/B _09288_/C vssd1 vssd1 vccd1 vccd1 _09290_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _11320_/A _11320_/B vssd1 vssd1 vccd1 vccd1 _11320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08305__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ _11250_/B _11250_/C _11250_/A vssd1 vssd1 vccd1 vccd1 _11252_/C sky130_fd_sc_hd__a21o_1
XANTENNA__10238__S1 _10429_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ _10199_/A _10200_/X _10046_/X _10050_/B vssd1 vssd1 vccd1 vccd1 _10202_/Y
+ sky130_fd_sc_hd__o211ai_2
X_11182_ _11371_/A _11180_/Y _10990_/B _10992_/B vssd1 vssd1 vccd1 vccd1 _11183_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11760__A0 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10133_ _11605_/A _10304_/C _10304_/D _11569_/A vssd1 vssd1 vccd1 vccd1 _10135_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10064_ _10065_/A _10065_/B _10065_/C vssd1 vssd1 vccd1 vccd1 _10064_/X sky130_fd_sc_hd__and3_1
X_14941_ _15214_/CLK _14941_/D vssd1 vssd1 vccd1 vccd1 _14941_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__10315__A1 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10315__B2 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14872_ _14876_/CLK _14872_/D vssd1 vssd1 vccd1 vccd1 _14872_/Q sky130_fd_sc_hd__dfxtp_1
X_13823_ _15383_/CLK hold762/X vssd1 vssd1 vccd1 vccd1 hold761/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10618__A2 _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13754_ _11104_/A _12261_/B _13753_/Y _07391_/Y vssd1 vssd1 vccd1 vccd1 _13754_/X
+ sky130_fd_sc_hd__a211o_1
X_10966_ _11597_/A _11573_/B _14966_/Q _11596_/A vssd1 vssd1 vccd1 vccd1 _10969_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12705_ _13080_/A1 _12704_/X _12702_/X vssd1 vssd1 vccd1 vccd1 _13155_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__13017__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13685_ hold1275/X _13718_/A1 _13698_/S vssd1 vssd1 vccd1 vccd1 _13685_/X sky130_fd_sc_hd__mux2_1
X_10897_ _11038_/B _10894_/Y _10669_/Y _10673_/C vssd1 vssd1 vccd1 vccd1 _10897_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08119__S0 _08130_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10448__C _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15424_ _15424_/CLK _15424_/D vssd1 vssd1 vccd1 vccd1 _15424_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12636_ _12642_/A1 _12635_/X _12700_/S0 vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_183_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ _15356_/CLK _15355_/D vssd1 vssd1 vccd1 vccd1 _15355_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11043__A2 _15223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12240__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _12692_/A1 _12566_/X _12366_/A vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08995__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306_ _15435_/CLK _14306_/D vssd1 vssd1 vccd1 vccd1 _14306_/Q sky130_fd_sc_hd__dfxtp_1
X_11518_ _11518_/A _11518_/B vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15286_ _15383_/CLK _15286_/D vssd1 vssd1 vccd1 vccd1 _15286_/Q sky130_fd_sc_hd__dfxtp_1
X_12498_ hold179/A hold345/A _14596_/Q _13965_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12498_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_123_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ _15434_/CLK _14237_/D vssd1 vssd1 vccd1 vccd1 _14237_/Q sky130_fd_sc_hd__dfxtp_1
X_11449_ _11449_/A _11449_/B _11607_/A _11448_/X vssd1 vssd1 vccd1 vccd1 _11607_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10183__C _10830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09095__S1 _10087_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ _15453_/CLK hold358/X vssd1 vssd1 vccd1 vccd1 hold357/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13129_/A hold67/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__and2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14105_/CLK hold146/X vssd1 vssd1 vccd1 vccd1 _14099_/Q sky130_fd_sc_hd__dfxtp_1
X_06990_ _13662_/A1 hold2071/X _06994_/S vssd1 vssd1 vccd1 vccd1 _06990_/X sky130_fd_sc_hd__mux2_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09172__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ _08989_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _08660_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07611_ hold2029/X _12329_/A _07626_/S vssd1 vssd1 vccd1 vccd1 _07611_/X sky130_fd_sc_hd__mux2_1
X_08591_ _08591_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08592_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ hold825/X _13746_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold826/A sky130_fd_sc_hd__mux2_1
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10639__B _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold2772_A _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07473_ hold243/X _07473_/B vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__and2_1
XANTENNA__13730__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ hold2331/X _09344_/B _09346_/B vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09143_ _09143_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ hold2762/X _09073_/Y _12256_/A vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08125__A _08869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12519__C1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08025_ _08526_/B _12221_/B vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout2 fanout2/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__buf_4
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11189__C _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 hold720/A vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold731 hold731/A vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold742 hold742/A vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold753 hold753/A vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 hold764/A vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold775 hold775/A vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_A _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 hold797/A vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _10183_/A _09979_/B _09676_/D _09979_/C _09828_/X vssd1 vssd1 vccd1 vccd1
+ _09984_/A sky130_fd_sc_hd__a41o_1
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2110 _11662_/X vssd1 vssd1 vccd1 vccd1 _14465_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2121 _15266_/Q vssd1 vssd1 vccd1 vccd1 hold2121/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07175__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2132 _13659_/X vssd1 vssd1 vccd1 vccd1 _15366_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08927_ _10700_/A _09712_/A _08926_/C _09039_/A vssd1 vssd1 vccd1 vccd1 _08928_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2143 _14356_/Q vssd1 vssd1 vccd1 vccd1 hold2143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_A _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2154 _07069_/X vssd1 vssd1 vccd1 vccd1 _13885_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2165 _14224_/Q vssd1 vssd1 vccd1 vccd1 hold2165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1420 _07634_/X vssd1 vssd1 vccd1 vccd1 _14257_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2176 _07049_/X vssd1 vssd1 vccd1 vccd1 _13865_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 _14669_/Q vssd1 vssd1 vccd1 vccd1 hold1431/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1442 _07641_/X vssd1 vssd1 vccd1 vccd1 _14264_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2187 _13897_/Q vssd1 vssd1 vccd1 vccd1 hold2187/X sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ _15146_/Q _09925_/A2 _13570_/B vssd1 vssd1 vccd1 vccd1 _08858_/Y sky130_fd_sc_hd__a21oi_1
Xhold2198 _11897_/X vssd1 vssd1 vccd1 vccd1 _14718_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _14115_/Q vssd1 vssd1 vccd1 vccd1 hold1453/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1464 _07742_/X vssd1 vssd1 vccd1 vccd1 _14361_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1475 _14131_/Q vssd1 vssd1 vccd1 vccd1 hold1475/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1486 _07582_/X vssd1 vssd1 vccd1 vccd1 _14206_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07809_ hold473/X _13714_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _15428_/Q vssd1 vssd1 vccd1 vccd1 hold1497/X sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ _08692_/A _08691_/B _08691_/A vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__o21ba_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ _10819_/B _10819_/C _10819_/A vssd1 vssd1 vccd1 vccd1 _10856_/B sky130_fd_sc_hd__a21o_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09403__B _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__A _14995_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10751_ _13588_/A _10751_/B vssd1 vssd1 vccd1 vccd1 _11113_/C sky130_fd_sc_hd__and2_1
XFILLER_0_211_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _13501_/A hold245/X vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__and2_1
X_10682_ _10681_/A _10681_/B _10681_/C vssd1 vssd1 vccd1 vccd1 _10684_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ hold949/A _15265_/Q _15073_/Q _14366_/Q _12459_/S _12474_/S1 vssd1 vssd1
+ vccd1 vccd1 _12421_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12222__A1 _12221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08977__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15140_ _15305_/CLK _15140_/D vssd1 vssd1 vccd1 vccd1 _15140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12352_ _12700_/S1 _12341_/X _12345_/X _12351_/X vssd1 vssd1 vccd1 vccd1 _12352_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _11497_/A _11302_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _11303_/X sky130_fd_sc_hd__o21a_1
X_15071_ _15360_/CLK _15071_/D vssd1 vssd1 vccd1 vccd1 _15071_/Q sky130_fd_sc_hd__dfxtp_1
X_12283_ _13171_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _14932_/D sky130_fd_sc_hd__nor2_2
X_14022_ _15460_/CLK _14022_/D vssd1 vssd1 vccd1 vccd1 _14022_/Q sky130_fd_sc_hd__dfxtp_1
X_11234_ _11234_/A _11234_/B vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11165_ _11605_/A _11606_/B _11570_/B _11569_/A vssd1 vssd1 vccd1 vccd1 _11165_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07085__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__A2 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _10115_/B _14959_/Q _10115_/D _10115_/A vssd1 vssd1 vccd1 vccd1 _10117_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12908__S0 _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11096_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11096_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10047_ _10046_/B _10046_/C _10046_/A vssd1 vssd1 vccd1 vccd1 _10047_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14924_ _15244_/CLK _14924_/D vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10839__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__C1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14855_ _15004_/CLK _14855_/D vssd1 vssd1 vccd1 vccd1 _14855_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13806_ _14783_/CLK _13806_/D vssd1 vssd1 vccd1 vccd1 _13806_/Q sky130_fd_sc_hd__dfxtp_1
X_14786_ _15440_/CLK _14786_/D vssd1 vssd1 vccd1 vccd1 _14786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ _14094_/Q _12126_/C vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__or2_2
XANTENNA__10459__B _11588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13737_ hold915/X _13737_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold916/A sky130_fd_sc_hd__mux2_1
XFILLER_0_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10949_ hold2781/X input21/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13200_/B sky130_fd_sc_hd__mux2_2
XANTENNA__12461__A1 _12642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _14971_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13668_ hold373/X _13668_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold374/A sky130_fd_sc_hd__mux2_1
XFILLER_0_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15444_/CLK _15407_/D vssd1 vssd1 vccd1 vccd1 _15407_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11016__A2 _11537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ _12700_/S0 _12614_/X _12618_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12620_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ _11645_/B _11650_/B _13598_/X _13459_/A vssd1 vssd1 vccd1 vccd1 _15325_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10224__B1 _11640_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ _15357_/CLK _15338_/D vssd1 vssd1 vccd1 vccd1 _15338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09090__B1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10775__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07640__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15269_ _15400_/CLK _15269_/D vssd1 vssd1 vccd1 vccd1 _15269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13713__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__A1 _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B2 _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2520_A _07389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _09827_/Y _09828_/X _09709_/D _09711_/A vssd1 vssd1 vccd1 vccd1 _09831_/C
+ sky130_fd_sc_hd__o211ai_2
Xfanout507 _06926_/Y vssd1 vssd1 vccd1 vccd1 _11303_/B1 sky130_fd_sc_hd__buf_8
Xfanout518 _15426_/Q vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__buf_8
XFILLER_0_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout529 _08869_/A vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__clkbuf_8
X_09761_ _09478_/A _09476_/X _09616_/A _09760_/Y _09759_/D vssd1 vssd1 vccd1 vccd1
+ _09763_/A sky130_fd_sc_hd__o311a_1
X_06973_ _14082_/Q _14091_/Q _06967_/X _11997_/B vssd1 vssd1 vccd1 vccd1 _06973_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08712_ _08712_/A _08712_/B _08712_/C vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__and3_2
XFILLER_0_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13725__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _09692_/A _09692_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09693_/A sky130_fd_sc_hd__and3_1
XFILLER_0_193_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07723__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08643_ hold2531/X _11643_/B _08256_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _08643_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08574_ _08893_/A _09008_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _08574_/X sky130_fd_sc_hd__and3_1
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12820__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ hold555/X hold2822/X _07528_/S vssd1 vssd1 vccd1 vccd1 hold556/A sky130_fd_sc_hd__mux2_1
XFILLER_0_194_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14840_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_A _07710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07456_ _07456_/A _13459_/A vssd1 vssd1 vccd1 vccd1 _14086_/D sky130_fd_sc_hd__and2_1
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12970__C_N _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A _15210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _14051_/Q _12308_/A _07387_/C _07387_/D vssd1 vssd1 vccd1 vccd1 _12379_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_0_88_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09126_ _10002_/C _09726_/B _09125_/C _09125_/D vssd1 vssd1 vccd1 vccd1 _09127_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_161_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09081__B1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ _09055_/B _09055_/C _09055_/A vssd1 vssd1 vccd1 vccd1 _09057_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ _08007_/B _08007_/C _08007_/A vssd1 vssd1 vccd1 vccd1 _08010_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__08005__D _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__A1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold550 hold550/A vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 hold561/A vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 hold572/A vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 hold583/A vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold594 hold594/A vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _10338_/B _11536_/B _10166_/C _10166_/A vssd1 vssd1 vccd1 vccd1 _09959_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _12970_/A _12970_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _12977_/B sky130_fd_sc_hd__or3b_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 _11841_/X vssd1 vssd1 vccd1 vccd1 _14664_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1261 _13815_/Q vssd1 vssd1 vccd1 vccd1 hold1261/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07633__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _11921_/A0 hold1897/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__mux2_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1272 _11684_/X vssd1 vssd1 vccd1 vccd1 _14487_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _15275_/Q vssd1 vssd1 vccd1 vccd1 hold1283/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1294 _07601_/X vssd1 vssd1 vccd1 vccd1 _14225_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08990__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14640_ _15444_/CLK _14640_/D vssd1 vssd1 vccd1 vccd1 _14640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ hold445/X _13739_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold446/A sky130_fd_sc_hd__mux2_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _11590_/A _11569_/B _11563_/B _11598_/A vssd1 vssd1 vccd1 vccd1 _10807_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11246__A2 _15221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12443__A1 _12474_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14571_ _15441_/CLK hold232/X vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__dfxtp_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ hold613/X _13703_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold614/A sky130_fd_sc_hd__mux2_1
XFILLER_0_200_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15357_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__A2 _13416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ _13736_/A1 hold1405/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13522_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _10734_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11651__C1 _13369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13453_ _10228_/B _13468_/A _13452_/Y _13797_/C1 vssd1 vssd1 vccd1 vccd1 _15220_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ _10664_/A _10664_/B _10664_/C vssd1 vssd1 vccd1 vccd1 _10666_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _13377_/B _12325_/B _12403_/X vssd1 vssd1 vccd1 vccd1 _12404_/X sky130_fd_sc_hd__a21o_1
X_13384_ _13389_/A _13384_/B vssd1 vssd1 vccd1 vccd1 _15175_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_152_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11954__A0 _13742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ _11320_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__nor2_1
X_15123_ _15132_/CLK _15123_/D vssd1 vssd1 vccd1 vccd1 _15123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12335_ _14331_/Q _14235_/Q _14395_/Q hold895/A _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12335_/X sky130_fd_sc_hd__mux4_1
XANTENNA__07808__S _07810_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15054_ _15278_/CLK _15054_/D vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__dfxtp_1
X_12266_ _13373_/A _13418_/B vssd1 vssd1 vccd1 vccd1 _14915_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_121_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _14409_/CLK hold714/X vssd1 vssd1 vccd1 vccd1 hold713/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09375__A1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _11370_/B _11215_/X _10994_/B _10996_/C vssd1 vssd1 vccd1 vccd1 _11217_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ hold165/A hold529/A _12198_/S vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_208_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08212__B _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11148_ _11578_/C _11148_/B _11148_/C vssd1 vssd1 vccd1 vccd1 _11434_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_208_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11079_ _11075_/Y _11077_/X _10852_/X _10856_/C vssd1 vssd1 vccd1 vccd1 _11080_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07543__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__B _11573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ _14992_/CLK _14907_/D vssd1 vssd1 vccd1 vccd1 _14907_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09043__B _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__D _08685_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14838_ _14842_/CLK _14838_/D vssd1 vssd1 vccd1 vccd1 _14838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14769_ _15411_/CLK _14769_/D vssd1 vssd1 vccd1 vccd1 _14769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk clkbuf_4_7__f_clk/X vssd1 vssd1 vccd1 vccd1 _15293_/CLK sky130_fd_sc_hd__clkbuf_16
X_07310_ _11378_/D _10283_/C vssd1 vssd1 vccd1 vccd1 _09619_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08290_ _08901_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__and2_1
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_9_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07241_ _10356_/C _10010_/B vssd1 vssd1 vccd1 vccd1 _07241_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15211__D _15211_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07172_ _13673_/A1 hold1663/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07718__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08403__A _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12596__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09813_ _09813_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09815_/B sky130_fd_sc_hd__nand2_1
Xfanout359 _12327_/A vssd1 vssd1 vccd1 vccd1 _13080_/A1 sky130_fd_sc_hd__buf_12
XANTENNA_fanout386_A _11762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09744_ _09745_/A _09745_/B _09745_/C _09745_/D vssd1 vssd1 vccd1 vccd1 _09744_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06956_ hold65/A hold321/A _06955_/X _14029_/Q vssd1 vssd1 vccd1 vccd1 _06956_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08776__C _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09234__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09675_ _09979_/B _09860_/B _09676_/D _10183_/A vssd1 vssd1 vccd1 vccd1 _09678_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout553_A _15423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__A2 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__D _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _08624_/X _08625_/Y _08515_/X _08517_/X vssd1 vssd1 vccd1 vccd1 _08629_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_A _14965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ _08981_/A _08557_/B vssd1 vssd1 vccd1 vccd1 _08557_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout818_A _14489_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _15077_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11703__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07508_ hold1907/X _13714_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07508_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ _08581_/B _08487_/C _08487_/A vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10827__B _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07439_ _07439_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14069_/D sky130_fd_sc_hd__nor2_1
XANTENNA__13203__B _13203_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12728__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ _11598_/A _11605_/B _10450_/C _10450_/D vssd1 vssd1 vccd1 vccd1 _10452_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11936__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09109_ _09514_/A _09109_/B vssd1 vssd1 vccd1 vccd1 _09109_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10381_ _10380_/A _10380_/B _10439_/B _10380_/D vssd1 vssd1 vccd1 vccd1 _10381_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12534__S _12560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ _12120_/A _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12120_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__07628__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12051_ _12059_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _14838_/D sky130_fd_sc_hd__and2_1
Xhold380 hold380/A vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold391 hold391/A vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ _11542_/B _11001_/X _11000_/X vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08565__C1 _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout860 _07473_/B vssd1 vssd1 vccd1 vccd1 _07474_/B sky130_fd_sc_hd__buf_4
XANTENNA__12339__S1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout871 _13486_/A vssd1 vssd1 vccd1 vccd1 _13487_/A sky130_fd_sc_hd__buf_2
XFILLER_0_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout882 _13381_/A vssd1 vssd1 vccd1 vccd1 _13373_/A sky130_fd_sc_hd__buf_4
Xfanout893 _13338_/A vssd1 vssd1 vccd1 vccd1 _13317_/A sky130_fd_sc_hd__buf_8
XFILLER_0_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _13742_/A1 _12329_/B _12953_/B1 _13197_/B vssd1 vssd1 vccd1 vccd1 _12953_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1080 _07807_/X vssd1 vssd1 vccd1 vccd1 _14422_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 _14395_/Q vssd1 vssd1 vccd1 vccd1 hold1091/X sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _13659_/A1 hold1051/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__mux2_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ hold329/A _13917_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__mux2_1
XANTENNA_220 _13444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08983__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10770__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _15045_/CLK hold764/X vssd1 vssd1 vccd1 vccd1 hold763/A sky130_fd_sc_hd__dfxtp_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11835_ hold435/X hold2783/X _11845_/S vssd1 vssd1 vccd1 vccd1 hold436/A sky130_fd_sc_hd__mux2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12709__S _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_clk clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 _14750_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14554_ _15456_/CLK _14554_/D vssd1 vssd1 vccd1 vccd1 _14554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ hold1401/X _13653_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11766_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _13653_/A1 hold1043/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13505_/X sky130_fd_sc_hd__mux2_1
X_10717_ _10717_/A _10717_/B _10717_/C vssd1 vssd1 vccd1 vccd1 _10719_/C sky130_fd_sc_hd__nand3_2
XANTENNA__07843__A1 _15342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08191__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14485_ _14485_/CLK _14485_/D vssd1 vssd1 vccd1 vccd1 _14485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11697_ hold289/X _13651_/A1 _11712_/S vssd1 vssd1 vccd1 vccd1 hold290/A sky130_fd_sc_hd__mux2_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10456__C _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ _09083_/A _12275_/B _13440_/S vssd1 vssd1 vccd1 vccd1 _13437_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_153_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10648_ _10473_/X _10476_/X _10646_/Y _10647_/X vssd1 vssd1 vccd1 vccd1 _10648_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11927__A0 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__A2 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13367_ _13369_/A _13367_/B vssd1 vssd1 vccd1 vccd1 _15158_/D sky130_fd_sc_hd__nor2_1
X_10579_ _11497_/A _10578_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _10579_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15106_ _15116_/CLK _15106_/D vssd1 vssd1 vccd1 vccd1 _15106_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07538__S _07544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12318_ hold589/A hold289/A hold855/A _14717_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12318_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_107_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13298_ input74/X fanout2/X _13297_/X vssd1 vssd1 vccd1 vccd1 _13299_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ _15427_/CLK _15037_/D vssd1 vssd1 vccd1 vccd1 _15037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12249_ _12243_/A _12248_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _12249_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2709 _12004_/X vssd1 vssd1 vccd1 vccd1 _12005_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07790_ hold781/X _13728_/A1 _07794_/S vssd1 vssd1 vccd1 vccd1 hold782/A sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12655__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09520__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _09599_/A _09459_/C _09459_/A vssd1 vssd1 vccd1 vccd1 _09461_/D sky130_fd_sc_hd__a21o_1
XANTENNA__12750__S1 _12944_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10761__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ _08411_/A _08468_/B _08411_/C vssd1 vssd1 vccd1 vccd1 _08474_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_203_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _09390_/A _09390_/B _09390_/C vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15296_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_176_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10607__A2_N _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A1 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _07900_/B _13382_/B _08287_/X vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13080__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07834__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ _12247_/A _08270_/X _08272_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _08274_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07224_ _12254_/A _07224_/B vssd1 vssd1 vccd1 vccd1 _07323_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07155_ _13656_/A1 hold2223/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07086_ _13689_/A1 hold2209/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07086_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09339__A1 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10497__B1_N _10482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12894__A1 _13050_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A _10700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ _14785_/Q hold483/A hold521/A _14721_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07989_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07183__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ _09727_/A _09727_/B vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__or2_1
X_06939_ _06939_/A vssd1 vssd1 vccd1 vccd1 _06939_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12102__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _10338_/B _09979_/D _09809_/C _10166_/A vssd1 vssd1 vccd1 vccd1 _09661_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08609_ _08610_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_194_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A _09589_/B vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__xnor2_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11620_ _11620_/A _11620_/B vssd1 vssd1 vccd1 vccd1 _11621_/B sky130_fd_sc_hd__nand2_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ _11551_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _11552_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07825__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ _10502_/A _10502_/B _10502_/C _10502_/D vssd1 vssd1 vccd1 vccd1 _10502_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14270_ _15434_/CLK _14270_/D vssd1 vssd1 vccd1 vccd1 _14270_/Q sky130_fd_sc_hd__dfxtp_1
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13221_ hold943/X _13519_/A0 _13236_/S vssd1 vssd1 vccd1 vccd1 hold944/A sky130_fd_sc_hd__mux2_1
X_10433_ _10433_/A _10433_/B vssd1 vssd1 vccd1 vccd1 _10433_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13152_ _13389_/A _13152_/B vssd1 vssd1 vccd1 vccd1 _15017_/D sky130_fd_sc_hd__nor2_1
X_10364_ _10364_/A _10364_/B _10364_/C vssd1 vssd1 vccd1 vccd1 _10364_/X sky130_fd_sc_hd__and3_2
XFILLER_0_131_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ hold2408/X _12129_/A2 _12102_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12103_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ hold1255/X hold1641/X hold571/X hold1389/X _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13083_/X sky130_fd_sc_hd__mux4_1
X_10295_ _10296_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10295_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11137__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ hold2439/X hold2678/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11688__A2 _13792_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07987__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07093__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 _13698_/A1 vssd1 vssd1 vccd1 vccd1 _13665_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12637__A1 _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13985_ _15385_/CLK _13985_/D vssd1 vssd1 vccd1 vccd1 _13985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__A1 _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _13092_/A1 _12935_/X _13050_/S0 vssd1 vssd1 vccd1 vccd1 _12936_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07821__S _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8__f_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12867_ _06942_/Y _12866_/X _14490_/Q vssd1 vssd1 vccd1 vccd1 _12867_/X sky130_fd_sc_hd__a21o_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ hold323/X _15058_/Q _11828_/S vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__mux2_1
X_14606_ _15373_/CLK _14606_/D vssd1 vssd1 vccd1 vccd1 _14606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12496__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12798_ hold217/A hold537/A hold613/A _13977_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12798_/X sky130_fd_sc_hd__mux4_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14537_ _15440_/CLK _14537_/D vssd1 vssd1 vccd1 vccd1 _14537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ _13735_/A1 hold1067/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11749_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14468_ _14731_/CLK _14468_/D vssd1 vssd1 vccd1 vccd1 _14468_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12248__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13419_ _08179_/B _13466_/A _13418_/Y _13178_/A vssd1 vssd1 vccd1 vccd1 _15203_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12799__S1 _12899_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _15391_/CLK _14399_/D vssd1 vssd1 vccd1 vccd1 _14399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10584__C1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08792__A2 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08960_ _07230_/A _07327_/B _08845_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _08960_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15301_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07911_ _07904_/A _07904_/B _07429_/A vssd1 vssd1 vccd1 vccd1 _07911_/X sky130_fd_sc_hd__a21o_1
Xhold2506 _15322_/Q vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08891_ _09008_/A _09864_/C _09864_/D _08893_/A vssd1 vssd1 vccd1 vccd1 _08895_/C
+ sky130_fd_sc_hd__a22o_1
Xhold2517 _08176_/Y vssd1 vssd1 vccd1 vccd1 _13418_/B sky130_fd_sc_hd__buf_1
XFILLER_0_209_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2528 _11649_/X vssd1 vssd1 vccd1 vccd1 hold2528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2539 _12159_/X vssd1 vssd1 vccd1 vccd1 _14890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1805 _13931_/Q vssd1 vssd1 vccd1 vccd1 hold1805/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07842_ _07862_/C _14031_/Q _14035_/Q _06908_/Y _07839_/X vssd1 vssd1 vccd1 vccd1
+ _07842_/X sky130_fd_sc_hd__o221a_1
Xhold1816 _07136_/X vssd1 vssd1 vccd1 vccd1 _13946_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1827 _14146_/Q vssd1 vssd1 vccd1 vccd1 hold1827/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12971__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08400__B _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1838 _07671_/X vssd1 vssd1 vccd1 vccd1 _14292_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1849 _13894_/Q vssd1 vssd1 vccd1 vccd1 hold1849/X sky130_fd_sc_hd__dlygate4sd3_1
X_07773_ _13744_/A1 hold1967/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07773_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__B2 _13184_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13733__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _09514_/A _09512_/B vssd1 vssd1 vccd1 vccd1 _09512_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12723__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07731__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09443_ _10110_/A _09724_/C _09724_/D _10002_/C vssd1 vssd1 vccd1 vccd1 _09445_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09512__A _09514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _10244_/A _09373_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _09374_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13053__A1 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13053__B2 _13201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08325_ _08324_/B _08324_/C _08324_/A vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout516_A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ _08256_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _08261_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_172_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09104__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07207_ hold1135/X _13741_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 _07207_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08187_ hold179/A hold345/A _14596_/Q _13965_/Q _08548_/S0 _08548_/S1 vssd1 vssd1
+ vccd1 vccd1 _08187_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_81_clk_A clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__S _07181_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07138_ _13739_/A1 hold1299/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07138_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09980__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__B _11614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07069_ _13674_/A1 hold2153/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07069_/X sky130_fd_sc_hd__mux2_1
Xoutput260 _14877_/Q vssd1 vssd1 vccd1 vccd1 out0[0] sky130_fd_sc_hd__buf_12
Xoutput271 _14878_/Q vssd1 vssd1 vccd1 vccd1 out0[1] sky130_fd_sc_hd__buf_12
Xoutput282 _14879_/Q vssd1 vssd1 vccd1 vccd1 out0[2] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12867__A1 _06942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _11288_/A1 _13396_/B _09956_/X vssd1 vssd1 vccd1 vccd1 _13450_/B sky130_fd_sc_hd__a21oi_4
XANTENNA_clkbuf_leaf_96_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput293 _14855_/Q vssd1 vssd1 vccd1 vccd1 out1[10] sky130_fd_sc_hd__buf_12
XANTENNA__10840__B _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12619__A1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12714__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ hold231/X vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__13292__A1 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _11605_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07641__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12721_ hold767/A _15277_/Q hold943/A _14378_/Q _12791_/S _12749_/S1 vssd1 vssd1
+ vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_179_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_154_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10568__A _10744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15440_ _15440_/CLK _15440_/D vssd1 vssd1 vccd1 vccd1 _15440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ _13027_/A _12652_/B _12652_/C vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__and3_1
XFILLER_0_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13044__A1 _13100_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _11603_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__xnor2_1
X_15371_ _15371_/CLK hold460/X vssd1 vssd1 vccd1 vccd1 hold459/A sky130_fd_sc_hd__dfxtp_1
X_12583_ hold777/A _14536_/Q _14696_/Q _14760_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12583_/X sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_169_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14322_ _15090_/CLK hold298/X vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11534_ _11341_/A _11341_/B _11338_/X vssd1 vssd1 vccd1 vccd1 _11535_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__08471__A1 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13598__B _13634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14253_ _15449_/CLK _14253_/D vssd1 vssd1 vccd1 vccd1 _14253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _11465_/A _11465_/B _11465_/C vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_leaf_49_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08759__C1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09646__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ _13716_/A _13650_/B vssd1 vssd1 vccd1 vccd1 _13204_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _10252_/A _10415_/X _11303_/B1 vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__o21a_1
X_14184_ _15184_/CLK hold144/X vssd1 vssd1 vccd1 vccd1 _14184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _11209_/A _11209_/C _11209_/B vssd1 vssd1 vccd1 vccd1 _11397_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__12650__S0 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output170_A _15182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ _13499_/A hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__and2_1
X_10347_ _10347_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10350_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07816__S _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ hold657/A _14264_/Q _13066_/S vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__mux2_1
X_10278_ _11597_/A _14961_/Q vssd1 vssd1 vccd1 vccd1 _10279_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _12059_/A _12017_/B vssd1 vssd1 vccd1 vccd1 _14821_/D sky130_fd_sc_hd__and2_1
XANTENNA__09723__B2 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08220__B _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _15400_/CLK _13968_/D vssd1 vssd1 vccd1 vccd1 _13968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _12950_/S0 _12914_/X _12918_/X _12944_/C1 vssd1 vssd1 vccd1 vccd1 _12920_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13899_ _15432_/CLK _13899_/D vssd1 vssd1 vccd1 vccd1 _13899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11801__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ hold2639/X _09925_/A2 _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08110_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ _15148_/Q _09925_/A2 _13570_/B vssd1 vssd1 vccd1 vccd1 _09090_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08462__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold2550_A _14829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08041_ _08256_/A _13346_/B vssd1 vssd1 vccd1 vccd1 _08046_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11349__A1 _11620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11349__B2 _11564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__S1 _09795_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 hold902/A vssd1 vssd1 vccd1 vccd1 hold902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold913 hold913/A vssd1 vssd1 vccd1 vccd1 hold913/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 hold924/A vssd1 vssd1 vccd1 vccd1 hold924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 hold935/A vssd1 vssd1 vccd1 vccd1 hold935/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__A1 _10022_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold946 hold946/A vssd1 vssd1 vccd1 vccd1 hold946/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13728__S _13732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold957 hold957/A vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__B2 _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold968 hold968/A vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _09989_/X _09990_/Y _09833_/X _09835_/Y vssd1 vssd1 vccd1 vccd1 _09993_/C
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__10941__A _11504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold979 hold979/A vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07726__S _07726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ _08939_/X _08941_/Y _08825_/B _08825_/Y vssd1 vssd1 vccd1 vccd1 _08944_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_110_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2303 _15293_/Q vssd1 vssd1 vccd1 vccd1 _07393_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07953__C _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2314 _14057_/Q vssd1 vssd1 vccd1 vccd1 _07852_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2325 _14918_/Q vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2336 hold2841/X vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__buf_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ hold799/A _14216_/Q hold701/A _14470_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08875_/B sky130_fd_sc_hd__mux4_1
Xhold2347 _13567_/X vssd1 vssd1 vccd1 vccd1 _15309_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 _13679_/X vssd1 vssd1 vccd1 vccd1 _15386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 _13971_/Q vssd1 vssd1 vccd1 vccd1 hold1613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2358 _10927_/X vssd1 vssd1 vccd1 vccd1 hold2358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2369 hold2837/X vssd1 vssd1 vccd1 vccd1 _08741_/A sky130_fd_sc_hd__buf_1
Xhold1624 _11669_/X vssd1 vssd1 vccd1 vccd1 _14472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1635 _14731_/Q vssd1 vssd1 vccd1 vccd1 hold1635/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 _07524_/X vssd1 vssd1 vccd1 vccd1 _14149_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07825_ _12247_/A _07820_/X _07824_/X _06926_/A vssd1 vssd1 vccd1 vccd1 _07826_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__D _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1657 _13856_/Q vssd1 vssd1 vccd1 vccd1 hold1657/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07820__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1668 _07099_/X vssd1 vssd1 vccd1 vccd1 _13912_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1679 _14143_/Q vssd1 vssd1 vccd1 vccd1 hold1679/X sky130_fd_sc_hd__dlygate4sd3_1
X_07756_ _13661_/A1 hold2139/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07756_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10088__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09810__A1_N _09661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07687_ hold1691/X _13512_/A0 _07693_/S vssd1 vssd1 vccd1 vccd1 _07687_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout633_A _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ _10000_/A _09846_/B _10283_/C vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__and3_1
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08128__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _09495_/A _09498_/C vssd1 vssd1 vccd1 vccd1 _09357_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout800_A _12689_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11711__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__S0 _11506_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _08222_/A _08222_/C _08222_/B vssd1 vssd1 vccd1 vccd1 _08310_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__08453__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _09288_/A _09288_/B _09288_/C vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__and3_1
XFILLER_0_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ _08239_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__A _14994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__B _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11250_ _11250_/A _11250_/B _11250_/C vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__nand3_2
XANTENNA__09402__B1 _15209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08205__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _10046_/X _10050_/B _10199_/A _10200_/X vssd1 vssd1 vccd1 vccd1 _10201_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11181_ _10990_/B _10992_/B _11371_/A _11180_/Y vssd1 vssd1 vccd1 vccd1 _11371_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__09953__B2 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07636__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _11569_/A _11605_/A _10304_/C _10304_/D vssd1 vssd1 vccd1 vccd1 _10135_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10063_ _10060_/Y _10061_/X _09898_/Y _09900_/Y vssd1 vssd1 vccd1 vccd1 _10065_/C
+ sky130_fd_sc_hd__a211o_1
X_14940_ _15292_/CLK _14940_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08064__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10315__A2 _14956_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ _14876_/CLK _14871_/D vssd1 vssd1 vccd1 vccd1 _14871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _15093_/CLK _13822_/D vssd1 vssd1 vccd1 vccd1 _13822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12699__S0 _12591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__A1 _06940_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13753_ _15134_/Q _07812_/A _13750_/A _13343_/B vssd1 vssd1 vccd1 vccd1 _13753_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
X_10965_ _11597_/A _11594_/B _10783_/X _10784_/X _11573_/B vssd1 vssd1 vccd1 vccd1
+ _10972_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12704_ _09079_/Y _13104_/A2 _12703_/X vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13017__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13684_ hold1767/X _15037_/Q _13698_/S vssd1 vssd1 vccd1 vccd1 _13684_/X sky130_fd_sc_hd__mux2_1
X_10896_ _10896_/A vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__inv_2
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08119__S1 _08130_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10448__D _11563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15423_ _15423_/CLK _15423_/D vssd1 vssd1 vccd1 vccd1 _15423_/Q sky130_fd_sc_hd__dfxtp_4
X_12635_ hold597/A _13939_/Q _12641_/S vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11123__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13402__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15354_ _15354_/CLK _15354_/D vssd1 vssd1 vccd1 vccd1 _15354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ hold319/A hold831/A _12566_/S vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12871__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ _11517_/A _15223_/Q vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14305_ _15264_/CLK hold346/X vssd1 vssd1 vccd1 vccd1 hold345/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15285_ _15382_/CLK hold626/X vssd1 vssd1 vccd1 vccd1 hold625/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12497_ _14788_/Q _14500_/Q _14628_/Q _14724_/Q _12460_/S _12689_/S1 vssd1 vssd1
+ vccd1 vccd1 _12497_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12528__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14236_ _15392_/CLK hold328/X vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__dfxtp_1
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ _11593_/B _11447_/C _11447_/A vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12623__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10183__D _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _14485_/CLK hold826/X vssd1 vssd1 vccd1 vccd1 hold825/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11379_ _11379_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11381_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13492_/A hold81/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__and2_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _15293_/CLK hold112/X vssd1 vssd1 vccd1 vccd1 _14098_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13891_/Q _14019_/Q hold945/A _13827_/Q _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13049_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08055__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09172__A2 _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07610_ _11730_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07610_/Y sky130_fd_sc_hd__nor2_4
X_08590_ _08589_/A _08589_/B _08589_/C vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__a21oi_1
X_07541_ hold493/X _13745_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold494/A sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2598_A _14427_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07472_ hold221/X _07474_/B vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ _09084_/B _09086_/B _09082_/X vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_17_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12767__B1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ _09140_/X _09142_/B vssd1 vssd1 vccd1 vccd1 _09143_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07310__A _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ _09119_/B _09073_/B vssd1 vssd1 vccd1 vccd1 _09073_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08024_ _08022_/Y _08024_/B vssd1 vssd1 vccd1 vccd1 _08024_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold710 hold710/A vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout3 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout3/X sky130_fd_sc_hd__buf_4
XFILLER_0_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12614__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold721 hold721/A vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 hold732/A vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__A2 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13458__S _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold743 hold743/A vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold754 hold754/A vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold765 hold765/A vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 hold776/A vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 hold787/A vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09975_ _09872_/A _09871_/B _09871_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__o21bai_2
Xhold798 hold798/A vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08141__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2100 _11706_/X vssd1 vssd1 vccd1 vccd1 _14502_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2111 _15071_/Q vssd1 vssd1 vccd1 vccd1 hold2111/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ _08926_/A _09712_/A _08926_/C _09039_/A vssd1 vssd1 vccd1 vccd1 _09039_/B
+ sky130_fd_sc_hd__nand4_2
Xhold2122 _13508_/X vssd1 vssd1 vccd1 vccd1 _15266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2133 _13933_/Q vssd1 vssd1 vccd1 vccd1 hold2133/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__B1 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2144 _07737_/X vssd1 vssd1 vccd1 vccd1 _14356_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1410 _07010_/X vssd1 vssd1 vccd1 vccd1 _13829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2155 _14331_/Q vssd1 vssd1 vccd1 vccd1 hold2155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2166 _07600_/X vssd1 vssd1 vccd1 vccd1 _14224_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1421 _13872_/Q vssd1 vssd1 vccd1 vccd1 hold1421/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2177 _14536_/Q vssd1 vssd1 vccd1 vccd1 hold2177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 _11846_/X vssd1 vssd1 vccd1 vccd1 _14669_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ _10233_/A _08857_/B _09087_/C vssd1 vssd1 vccd1 vccd1 _08857_/X sky130_fd_sc_hd__or3_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1443 _14006_/Q vssd1 vssd1 vccd1 vccd1 hold1443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2188 _07084_/X vssd1 vssd1 vccd1 vccd1 _13897_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1454 _07487_/X vssd1 vssd1 vccd1 vccd1 _14115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2199 _14554_/Q vssd1 vssd1 vccd1 vccd1 hold2199/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1465 _14233_/Q vssd1 vssd1 vccd1 vccd1 hold1465/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout848_A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__B1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ hold489/X _13746_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold490/A sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1476 _07503_/X vssd1 vssd1 vccd1 vccd1 _14131_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13247__A1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08788_ _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__xnor2_2
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1487 _14548_/Q vssd1 vssd1 vccd1 vccd1 hold1487/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07191__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1498 _13718_/X vssd1 vssd1 vccd1 vccd1 _15428_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ hold1095/X _13745_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07739_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09403__C _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12110__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11007__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10750_ _13750_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _10750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09409_ _09408_/B _09408_/C _09408_/A vssd1 vssd1 vccd1 vccd1 _09411_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12207__C1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _10681_/A _10681_/B _10681_/C vssd1 vssd1 vccd1 vccd1 _10684_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ _12420_/A _12420_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_106_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09623__B1 _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7__f_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7__f_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _12669_/A1 _12346_/X _12350_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_180_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _13892_/Q hold401/A _13860_/Q _13828_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _11302_/X sky130_fd_sc_hd__mux4_1
X_15070_ _15428_/CLK _15070_/D vssd1 vssd1 vccd1 vccd1 _15070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12282_ _13168_/A _13450_/B vssd1 vssd1 vccd1 vccd1 _14931_/D sky130_fd_sc_hd__nor2_2
X_14021_ _15387_/CLK _14021_/D vssd1 vssd1 vccd1 vccd1 _14021_/Q sky130_fd_sc_hd__dfxtp_1
X_11233_ _11340_/A _15225_/Q _11234_/A vssd1 vssd1 vccd1 vccd1 _11343_/B sky130_fd_sc_hd__and3_1
XFILLER_0_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _10972_/A _10972_/C _10972_/B vssd1 vssd1 vccd1 vccd1 _11179_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10115_ _10115_/A _10115_/B _14959_/Q _10115_/D vssd1 vssd1 vccd1 vccd1 _10115_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__12908__S1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11278_/B sky130_fd_sc_hd__and2_1
XANTENNA__07890__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ _10046_/A _10046_/B _10046_/C vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__or3_4
X_14923_ _15243_/CLK _14923_/D vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12694__C1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _15004_/CLK _14854_/D vssd1 vssd1 vccd1 vccd1 _14854_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _14397_/CLK hold746/X vssd1 vssd1 vccd1 vccd1 hold745/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11997_ _11997_/A _11997_/B _11997_/C _11997_/D vssd1 vssd1 vccd1 vccd1 _12128_/C
+ sky130_fd_sc_hd__or4_4
X_14785_ _15397_/CLK _14785_/D vssd1 vssd1 vccd1 vccd1 _14785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08665__A1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13736_ hold511/X _13736_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold512/A sky130_fd_sc_hd__mux2_1
X_10948_ _11320_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10879_ _11541_/A _11351_/B _11564_/B _11614_/B vssd1 vssd1 vccd1 vccd1 _10881_/C
+ sky130_fd_sc_hd__nand4_1
X_13667_ hold767/X _13700_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold768/A sky130_fd_sc_hd__mux2_1
XFILLER_0_27_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13097__S0 _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15443_/CLK hold406/X vssd1 vssd1 vccd1 vccd1 hold405/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ _12674_/S1 _12615_/X _12617_/X vssd1 vssd1 vccd1 vccd1 _12618_/X sky130_fd_sc_hd__a21o_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _13598_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13598_/X sky130_fd_sc_hd__or2_1
XANTENNA__13410__A1 _12262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15337_ _15340_/CLK _15337_/D vssd1 vssd1 vccd1 vccd1 _15337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ _13871_/Q _13999_/Q _13839_/Q _13807_/Q _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12549_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_1 _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _15268_/CLK _15268_/D vssd1 vssd1 vccd1 vccd1 _15268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09917__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14219_ _15276_/CLK _14219_/D vssd1 vssd1 vccd1 vccd1 _14219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15199_ _15199_/CLK _15199_/D vssd1 vssd1 vccd1 vccd1 _15199_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10527__A2 _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout508 _08065_/A vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__buf_6
Xfanout519 _15426_/Q vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__buf_6
XANTENNA__15209__D _15209_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ _09760_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09760_/Y sky130_fd_sc_hd__nand2_1
X_06972_ _14093_/Q _06972_/B _06972_/C _06972_/D vssd1 vssd1 vccd1 vccd1 _06972_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12910__S _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13021__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ _08805_/B _08709_/C _08709_/A vssd1 vssd1 vccd1 vccd1 _08712_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11488__B1 _13636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _09690_/B _09690_/C _09690_/A vssd1 vssd1 vccd1 vccd1 _09692_/C sky130_fd_sc_hd__a21o_1
X_08642_ _08642_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08573_ _09008_/A _09858_/A _09858_/B _08893_/A vssd1 vssd1 vccd1 vccd1 _08573_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13741__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07524_ hold1645/X _13728_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07524_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08200__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__A0 _13691_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07455_ _07455_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07455_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__A _10666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout429_A _11796_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07386_ _07438_/A _14060_/Q _07404_/A _15349_/Q _07385_/X vssd1 vssd1 vccd1 vccd1
+ _07387_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _10002_/C _09726_/B _09125_/C _09125_/D vssd1 vssd1 vccd1 vccd1 _09127_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_5_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11963__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _09056_/A vssd1 vssd1 vccd1 vccd1 _09056_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08007_ _08007_/A _08007_/B _08007_/C vssd1 vssd1 vccd1 vccd1 _08010_/B sky130_fd_sc_hd__or3_1
XFILLER_0_114_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout798_A _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold540 hold540/A vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08267__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold551 hold551/A vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__A2 _15220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 hold562/A vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07186__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold573 hold573/A vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold584 hold584/A vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold595 hold595/A vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_15__f_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_92_clk/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09958_ _09839_/B _09958_/B vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__nand2b_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _08909_/A _08909_/B _08909_/C vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__nand3_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09888_/B _09888_/C _09888_/A vssd1 vssd1 vccd1 vccd1 _09889_/X sky130_fd_sc_hd__a21o_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1240 _07507_/X vssd1 vssd1 vccd1 vccd1 _14135_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1251 _14289_/Q vssd1 vssd1 vccd1 vccd1 hold1251/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1262 _06996_/X vssd1 vssd1 vccd1 vccd1 _13815_/D sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ _13741_/A1 hold1241/X _11927_/S vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__mux2_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1273 _14279_/Q vssd1 vssd1 vccd1 vccd1 hold1273/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1284 _13517_/X vssd1 vssd1 vccd1 vccd1 _15275_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 _14258_/Q vssd1 vssd1 vccd1 vccd1 hold1295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ hold921/X _13738_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 hold922/A sky130_fd_sc_hd__mux2_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08990__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13651__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10802_ _10802_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10810_/A sky130_fd_sc_hd__nor2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14602_/CLK hold236/X vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__dfxtp_1
X_11782_ hold541/X _13669_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 hold542/A sky130_fd_sc_hd__mux2_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09430__A _10022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ _10733_/A _10733_/B vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__nand2_1
X_13521_ _13669_/A1 hold2169/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13521_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12795__C_N _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _13468_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13452_/Y sky130_fd_sc_hd__nand2_1
X_10664_ _10664_/A _10664_/B _10664_/C vssd1 vssd1 vccd1 vccd1 _10666_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_180_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ _13687_/A1 _12329_/B _12953_/B1 _13175_/B vssd1 vssd1 vccd1 vccd1 _12403_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ _13386_/A _13383_/B vssd1 vssd1 vccd1 vccd1 _15174_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _10580_/Y _10585_/Y _10594_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _10596_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15122_ _15132_/CLK _15122_/D vssd1 vssd1 vccd1 vccd1 _15122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _13373_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _14941_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15053_ _15278_/CLK _15053_/D vssd1 vssd1 vccd1 vccd1 _15053_/Q sky130_fd_sc_hd__dfxtp_1
X_12265_ _13150_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _14914_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_32_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07096__S _07096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ _14731_/CLK _14004_/D vssd1 vssd1 vccd1 vccd1 _14004_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12903__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ _10994_/B _10996_/C _11370_/B _11215_/X vssd1 vssd1 vccd1 vccd1 _11331_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output250_A _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ _13862_/Q _13990_/Q _13830_/Q _13798_/Q _12198_/S _12211_/S1 vssd1 vssd1
+ vccd1 vccd1 _12196_/X sky130_fd_sc_hd__mux4_1
XANTENNA_output348_A _14844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11147_ _11148_/B _11148_/C vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11078_ _10852_/X _10856_/C _11075_/Y _11077_/X vssd1 vssd1 vccd1 vccd1 _11080_/A
+ sky130_fd_sc_hd__a211oi_1
Xinput160 in2[9] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__clkbuf_2
X_10029_ _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1 _10044_/A sky130_fd_sc_hd__xnor2_2
X_14906_ _14992_/CLK _14906_/D vssd1 vssd1 vccd1 vccd1 _14906_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14837_ _14842_/CLK _14837_/D vssd1 vssd1 vccd1 vccd1 _14837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12419__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14768_ _15372_/CLK _14768_/D vssd1 vssd1 vccd1 vccd1 _14768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13719_ hold635/X _13719_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 hold636/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14699_ _15367_/CLK _14699_/D vssd1 vssd1 vccd1 vccd1 _14699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07240_ _07240_/A _07240_/B vssd1 vssd1 vccd1 vccd1 _11286_/A sky130_fd_sc_hd__and2_1
XFILLER_0_156_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07171_ _13705_/A1 hold1775/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07171_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold2728_A _15058_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08403__B _08776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13736__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ _09812_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__or2_1
XANTENNA__12640__S _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09743_ _09741_/A _09741_/B _09599_/B vssd1 vssd1 vccd1 vccd1 _09745_/D sky130_fd_sc_hd__o21ba_1
X_06955_ hold221/A hold257/A hold267/A hold243/A vssd1 vssd1 vccd1 vccd1 _06955_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout379_A _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ _10129_/A _11407_/A _09566_/X _09430_/X _09708_/B vssd1 vssd1 vccd1 vccd1
+ _09679_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08625_ _08621_/Y _08622_/X _08491_/A _08492_/B vssd1 vssd1 vccd1 vccd1 _08625_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A _13101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout546_A _15423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ hold631/A hold973/A hold781/A _14117_/Q _08990_/S0 _08990_/S1 vssd1 vssd1
+ vccd1 vccd1 _08557_/B sky130_fd_sc_hd__mux4_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07507_ hold1239/X _13680_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07507_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_194_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08487_ _08487_/A _08581_/B _08487_/C vssd1 vssd1 vccd1 vccd1 _08491_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10827__C _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07438_ _07438_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14068_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12808__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12189__A1 hold2564/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07369_ _07365_/X _07366_/Y _07367_/X _07368_/Y vssd1 vssd1 vccd1 vccd1 _07369_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12815__S _12915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13500__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ _14669_/Q _13942_/Q hold395/A _13910_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09109_/B sky130_fd_sc_hd__mux4_1
X_10380_ _10380_/A _10380_/B _10439_/B _10380_/D vssd1 vssd1 vccd1 vccd1 _10380_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__08262__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09039_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__A _14998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12050_ hold2555/X hold2720/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold370 hold370/A vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 hold381/A vssd1 vssd1 vccd1 vccd1 hold381/X sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _11586_/A _11614_/A _11378_/D vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__and3_1
Xhold392 hold392/A vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout850 _13455_/A vssd1 vssd1 vccd1 vccd1 _13477_/A sky130_fd_sc_hd__clkbuf_8
Xfanout861 _13455_/A vssd1 vssd1 vccd1 vccd1 _07473_/B sky130_fd_sc_hd__buf_2
Xfanout872 _13479_/A vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__buf_4
XFILLER_0_205_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout883 _13390_/A vssd1 vssd1 vccd1 vccd1 _13381_/A sky130_fd_sc_hd__clkbuf_8
Xfanout894 input161/X vssd1 vssd1 vccd1 vccd1 _13338_/A sky130_fd_sc_hd__buf_6
XFILLER_0_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12358__A2_N _08636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _13102_/A _12952_/B _12952_/C vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__and3_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 _11666_/X vssd1 vssd1 vccd1 vccd1 _14469_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1081 _14255_/Q vssd1 vssd1 vccd1 vccd1 hold1081/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _13691_/A1 hold1477/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11903_/X sky130_fd_sc_hd__mux2_1
Xhold1092 _07780_/X vssd1 vssd1 vccd1 vccd1 _14395_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12883_ hold679/A _14548_/Q hold325/A _14772_/Q _12941_/S _13024_/S1 vssd1 vssd1
+ vccd1 vccd1 _12883_/X sky130_fd_sc_hd__mux4_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07540__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_221 _13444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _15428_/CLK _14622_/D vssd1 vssd1 vccd1 vccd1 _14622_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10770__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11834_ hold1617/X _13721_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 _11834_/X sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ _15418_/CLK _14553_/D vssd1 vssd1 vccd1 vccd1 _14553_/Q sky130_fd_sc_hd__dfxtp_1
X_11765_ hold907/X _13652_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 hold908/A sky130_fd_sc_hd__mux2_1
XFILLER_0_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10716_ _10713_/Y _10714_/X _10498_/X _10502_/C vssd1 vssd1 vccd1 vccd1 _10717_/C
+ sky130_fd_sc_hd__o211ai_2
X_13504_ _13652_/A1 hold1355/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13504_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14484_ _14485_/CLK _14484_/D vssd1 vssd1 vccd1 vccd1 hold999/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11696_ _11730_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ _11564_/A _10827_/D _10646_/C _10646_/D vssd1 vssd1 vccd1 vccd1 _10647_/X
+ sky130_fd_sc_hd__a22o_1
X_13435_ _08966_/A _13440_/S _13434_/Y _13541_/A vssd1 vssd1 vccd1 vccd1 _15211_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13366_ _13369_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _15157_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10578_ _13888_/Q _14016_/Q _13856_/Q _13824_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _10578_/X sky130_fd_sc_hd__mux4_1
X_15105_ _15116_/CLK _15105_/D vssd1 vssd1 vccd1 vccd1 _15105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12317_ hold917/A _15261_/Q _15069_/Q _14362_/Q _12466_/S _12343_/A vssd1 vssd1 vccd1
+ vccd1 _12317_/X sky130_fd_sc_hd__mux4_1
X_13297_ input138/X fanout5/X fanout3/X input106/X vssd1 vssd1 vccd1 vccd1 _13297_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12248_ _15391_/Q _14526_/Q hold343/A _14750_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12248_/X sky130_fd_sc_hd__mux4_1
X_15036_ _15289_/CLK _15036_/D vssd1 vssd1 vccd1 vccd1 _15036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12888__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12352__A1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12460__S _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _12112_/A _12131_/X _12178_/X _13491_/A vssd1 vssd1 vccd1 vccd1 _12179_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08859__A1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07531__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _08503_/B _08410_/B vssd1 vssd1 vccd1 vccd1 _08411_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11804__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10761__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09390_ _09390_/A _09390_/B _09390_/C vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__and3_1
XANTENNA__09808__B1 _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08341_ hold2521/X _08526_/B _12221_/B _08340_/Y _08337_/Y vssd1 vssd1 vccd1 vccd1
+ _13382_/B sky130_fd_sc_hd__a221o_4
XFILLER_0_164_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08087__A2 _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold2678_A _14830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08272_ _08873_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08272_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07223_ _08677_/A _10873_/A vssd1 vssd1 vccd1 vccd1 _07224_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12635__S _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07047__A0 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12040__A0 hold2591/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07154_ _13655_/A1 hold1919/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07085_ _13721_/A1 hold1563/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07085_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13540__A0 _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07987_ hold949/A _15265_/Q _15073_/Q _14366_/Q _08130_/S0 _08130_/S1 vssd1 vssd1
+ vccd1 vccd1 _07987_/X sky130_fd_sc_hd__mux4_1
X_09726_ _10033_/A _09726_/B _09726_/C _09726_/D vssd1 vssd1 vccd1 vccd1 _09727_/B
+ sky130_fd_sc_hd__and4_1
X_06938_ _06938_/A vssd1 vssd1 vccd1 vccd1 _06938_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10657__A1 _11570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _09816_/A _10166_/C vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout830_A _12791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11714__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08608_ _08608_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__xor2_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09588_ _09589_/B _09589_/A vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__and2b_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08539_ _15143_/Q _09925_/A2 _09494_/A1 vssd1 vssd1 vccd1 vccd1 _08539_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_195_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11550_ _11550_/A _15224_/Q vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout6_A fanout6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ _10498_/X _10499_/Y _10323_/X _10328_/B vssd1 vssd1 vccd1 vccd1 _10502_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _11481_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__and2_1
XFILLER_0_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13220_ hold1259/X _13666_/A1 _13220_/S vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07639__S _07642_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10417_/Y _10422_/Y _10431_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _10433_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _13389_/A _13151_/B vssd1 vssd1 vccd1 vccd1 _15016_/D sky130_fd_sc_hd__nor2_1
X_10363_ _10362_/B _10362_/C _10362_/A vssd1 vssd1 vccd1 vccd1 _10364_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10593__B1 _11499_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _12102_/A _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12102_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13082_ _13107_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _14971_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_209_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10294_ _10294_/A _10294_/B vssd1 vssd1 vccd1 vccd1 _10296_/B sky130_fd_sc_hd__xor2_2
X_12033_ _12037_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _14829_/D sky130_fd_sc_hd__and2_1
XANTENNA__11685__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__B _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clk_A clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _13703_/A1 vssd1 vssd1 vccd1 vccd1 _13736_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout691 hold2823/X vssd1 vssd1 vccd1 vccd1 _13698_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08994__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ _15416_/CLK _13984_/D vssd1 vssd1 vccd1 vccd1 _13984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _14678_/Q _13951_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__mux2_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12866_ hold931/A hold699/A _12866_/S vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _15375_/CLK hold586/X vssd1 vssd1 vccd1 vccd1 hold585/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11817_ hold615/X _13671_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 hold616/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12496__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797_ hold455/A hold549/A _14640_/Q _14736_/Q _12735_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12797_/X sky130_fd_sc_hd__mux4_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _15042_/CLK _14536_/D vssd1 vssd1 vccd1 vccd1 _14536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11748_ _13734_/A1 hold693/X _11761_/S vssd1 vssd1 vccd1 vccd1 hold694/A sky130_fd_sc_hd__mux2_1
XFILLER_0_56_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14467_ _15080_/CLK _14467_/D vssd1 vssd1 vccd1 vccd1 _14467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12248__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _13743_/A1 hold2301/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12022__A0 _14984_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13140__A _13373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13418_ _13466_/A _13418_/B vssd1 vssd1 vccd1 vccd1 _13418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14398_ _15434_/CLK hold780/X vssd1 vssd1 vccd1 vccd1 hold779/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _13360_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _15140_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__S0 _11306_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07910_ _09344_/B _07910_/B vssd1 vssd1 vccd1 vccd1 _08964_/B sky130_fd_sc_hd__or2_2
XFILLER_0_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15019_ _15184_/CLK _15019_/D vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__dfxtp_1
X_08890_ _08890_/A _08890_/B vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_20_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2507 _13593_/X vssd1 vssd1 vccd1 vccd1 _15322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2518 _14874_/Q vssd1 vssd1 vccd1 vccd1 hold2518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2529 _14069_/Q vssd1 vssd1 vccd1 vccd1 _07411_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07841_ _14031_/Q _14032_/Q _07841_/C vssd1 vssd1 vccd1 vccd1 _07841_/X sky130_fd_sc_hd__or3_1
Xhold1806 _07121_/X vssd1 vssd1 vccd1 vccd1 _13931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1817 _13893_/Q vssd1 vssd1 vccd1 vccd1 hold1817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1828 _07521_/X vssd1 vssd1 vccd1 vccd1 _14146_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15217__D _15217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1839 _13871_/Q vssd1 vssd1 vccd1 vccd1 hold1839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_155_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07772_ hold2765/A hold1781/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07772_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12628__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09511_ _14285_/Q _14221_/Q hold417/A _14475_/Q _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09512_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10939__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B1 _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09454_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13038__C1 hold2774/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07313__A _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09373_ _15408_/Q _14543_/Q hold911/A hold863/A _10087_/S0 _10087_/S1 vssd1 vssd1
+ vccd1 vccd1 _09373_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13053__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08324_ _08324_/A _08324_/B _08324_/C vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__and3_1
XFILLER_0_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _13349_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout411_A _07080_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07206_ hold839/X _13674_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold840/A sky130_fd_sc_hd__mux2_1
XFILLER_0_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09104__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08186_ _13570_/B hold2688/X _08185_/X _13565_/C1 vssd1 vssd1 vccd1 vccd1 _08186_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08768__B1 _08992_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07137_ _13738_/A1 hold2089/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07137_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08863__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09980__A2 _11378_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__C _11378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _13673_/A1 hold1045/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07068_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout780_A _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput250 _14426_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[2] sky130_fd_sc_hd__buf_12
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout878_A _13479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput261 _14887_/Q vssd1 vssd1 vccd1 vccd1 out0[10] sky130_fd_sc_hd__buf_12
XANTENNA__11709__S _11712_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput272 _14897_/Q vssd1 vssd1 vccd1 vccd1 out0[20] sky130_fd_sc_hd__buf_12
Xoutput283 _14907_/Q vssd1 vssd1 vccd1 vccd1 out0[30] sky130_fd_sc_hd__buf_12
XANTENNA__10327__B1 _10326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput294 _14856_/Q vssd1 vssd1 vccd1 vccd1 out1[11] sky130_fd_sc_hd__buf_12
XFILLER_0_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07194__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09709_ _10129_/A _09709_/B _09709_/C _09709_/D vssd1 vssd1 vccd1 vccd1 _09711_/A
+ sky130_fd_sc_hd__nand4_2
X_10981_ _11606_/B _10980_/X _10979_/X vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__09496__A1 _13590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _12720_/A _12720_/B _13101_/A vssd1 vssd1 vccd1 vccd1 _12727_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07223__A _08677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12651_ _12676_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12652_/C sky130_fd_sc_hd__or2_1
XFILLER_0_167_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08038__B _08038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ _11602_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__xnor2_1
X_12582_ _12607_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _14951_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_26_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15370_ _15440_/CLK _15370_/D vssd1 vssd1 vccd1 vccd1 _15370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ _14612_/CLK hold336/X vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11533_ _11365_/A _11364_/B _11364_/A vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12004__A0 hold2548/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ _11465_/A _11465_/B _11465_/C vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__o21a_1
X_14252_ _15410_/CLK _14252_/D vssd1 vssd1 vccd1 vccd1 _14252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12555__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10415_ _13887_/Q _14015_/Q hold739/A hold761/A _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10415_/X sky130_fd_sc_hd__mux4_1
X_13203_ _13404_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _15068_/D sky130_fd_sc_hd__and2_1
XFILLER_0_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11395_ _11626_/A _11394_/C _11394_/A vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__a21o_1
X_14183_ _15184_/CLK hold150/X vssd1 vssd1 vccd1 vccd1 _14183_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08989__A _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12650__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _11340_/A _11620_/B vssd1 vssd1 vccd1 vccd1 _10347_/B sky130_fd_sc_hd__nand2_1
X_13134_ _13492_/A hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__and2_1
XANTENNA_output163_A _15175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13504__A0 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ hold473/X hold1907/X _13066_/S vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__mux2_1
X_10277_ _10275_/X _10277_/B vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12016_ hold2602/X hold2658/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12017_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09723__A2 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output330_A _14828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08220__C _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13967_ _15391_/CLK _13967_/D vssd1 vssd1 vccd1 vccd1 _13967_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13135__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ _12939_/S1 _12915_/X _12917_/X vssd1 vssd1 vccd1 vccd1 _12918_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_159_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13898_ _15433_/CLK _13898_/D vssd1 vssd1 vccd1 vccd1 _13898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12849_ _13883_/Q hold621/A hold397/A _13819_/Q _12915_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12849_/X sky130_fd_sc_hd__mux4_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08998__B1 _09724_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12794__A1 _12844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519_ _15063_/CLK hold684/X vssd1 vssd1 vccd1 vccd1 hold683/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08040_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _13346_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A2 _11614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 hold903/A vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 hold914/A vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold925 hold925/A vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 hold936/A vssd1 vssd1 vccd1 vccd1 hold936/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold947 hold947/A vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 hold958/A vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _09833_/X _09835_/Y _09989_/X _09990_/Y vssd1 vssd1 vccd1 vccd1 _09993_/B
+ sky130_fd_sc_hd__o211a_2
Xhold969 hold969/A vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2710_A _15165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _08825_/B _08825_/Y _08939_/X _08941_/Y vssd1 vssd1 vccd1 vccd1 _08944_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__12214__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__D _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2304 _07393_/X vssd1 vssd1 vccd1 vccd1 _14023_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2315 _14915_/Q vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold2326 _15311_/Q vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__buf_1
Xhold2337 _13543_/X vssd1 vssd1 vccd1 vccd1 _15297_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2348 _14060_/Q vssd1 vssd1 vccd1 vccd1 _06919_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08873_ _08873_/A _08873_/B vssd1 vssd1 vccd1 vccd1 _08873_/Y sky130_fd_sc_hd__nor2_1
Xhold1603 _14717_/Q vssd1 vssd1 vccd1 vccd1 hold1603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1614 _07163_/X vssd1 vssd1 vccd1 vccd1 _13971_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13744__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2359 _10928_/X vssd1 vssd1 vccd1 vccd1 _14451_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1625 _14134_/Q vssd1 vssd1 vccd1 vccd1 hold1625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1636 _11910_/X vssd1 vssd1 vccd1 vccd1 _14731_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07824_ _12233_/A _07821_/X _07823_/X vssd1 vssd1 vccd1 vccd1 _07824_/X sky130_fd_sc_hd__a21o_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1647 _13991_/Q vssd1 vssd1 vccd1 vccd1 hold1647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 _07039_/X vssd1 vssd1 vccd1 vccd1 _13856_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07820__S1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07742__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1669 _15430_/Q vssd1 vssd1 vccd1 vccd1 hold1669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09523__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ _13512_/A0 hold1121/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07755_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout361_A _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07686_ hold1131/X _13725_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 _07686_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09425_ _09846_/B _10010_/B _10283_/C _11580_/A vssd1 vssd1 vccd1 vccd1 _09457_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout626_A _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12234__B1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ _09350_/A _09222_/B _09355_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _09356_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10245__C1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__S1 _11506_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ _08306_/B _08306_/C _08306_/A vssd1 vssd1 vccd1 vccd1 _08310_/B sky130_fd_sc_hd__a21o_1
X_09287_ _09154_/A _09154_/B _09154_/C vssd1 vssd1 vccd1 vccd1 _09288_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__A1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10796__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07189__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ _08239_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12537__A1 _12668_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__C _09026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08169_ _07227_/B _08169_/B vssd1 vssd1 vccd1 vccd1 _08169_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09402__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10200_ _10198_/B _10198_/C _10198_/A vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ _11179_/B _11179_/C _11179_/A vssd1 vssd1 vccd1 vccd1 _11180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10131_ _11569_/A _11605_/A _10304_/C _10304_/D vssd1 vssd1 vccd1 vccd1 _10131_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12124__A _15002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12396__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10062_ _09898_/Y _09900_/Y _10060_/Y _10061_/X vssd1 vssd1 vccd1 vccd1 _10065_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__08064__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2860 _14067_/Q vssd1 vssd1 vccd1 vccd1 hold2860/X sky130_fd_sc_hd__dlygate4sd3_1
X_14870_ _14876_/CLK _14870_/D vssd1 vssd1 vccd1 vccd1 _14870_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07652__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ _14612_/CLK hold868/X vssd1 vssd1 vccd1 vccd1 hold867/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12699__S1 _12699_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__A2 _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _15459_/Q _07926_/A hold2366/X _13409_/A vssd1 vssd1 vccd1 vccd1 _13752_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10964_ _10964_/A _10964_/B vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ _13666_/A1 _13103_/A2 _13078_/B1 _13187_/B vssd1 vssd1 vccd1 vccd1 _12703_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13683_ _13683_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13715_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_211_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10895_ _10669_/Y _10673_/C _11038_/B _10894_/Y vssd1 vssd1 vccd1 vccd1 _10896_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_156_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11902__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15422_ _15422_/CLK _15422_/D vssd1 vssd1 vccd1 vccd1 _15422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12634_ _15440_/Q _13907_/Q _12641_/S vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12225__B1 _13172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12320__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11123__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15353_ _15354_/CLK _15353_/D vssd1 vssd1 vccd1 vccd1 _15353_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_109_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12565_ hold959/X hold561/X _12566_/S vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_182_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07099__S _07112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14304_ _14595_/CLK hold334/X vssd1 vssd1 vccd1 vccd1 hold333/A sky130_fd_sc_hd__dfxtp_1
X_11516_ _07264_/A _07287_/Y _11324_/X _11640_/B1 vssd1 vssd1 vccd1 vccd1 _11516_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15284_ _15408_/CLK _15284_/D vssd1 vssd1 vccd1 vccd1 _15284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ hold647/A _15268_/Q _15076_/Q _14369_/Q _12491_/S _12599_/S1 vssd1 vssd1
+ vccd1 vccd1 _12496_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12528__B2 _13180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14235_ _15360_/CLK _14235_/D vssd1 vssd1 vccd1 vccd1 _14235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _11447_/A _11593_/B _11447_/C vssd1 vssd1 vccd1 vccd1 _11607_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_46_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12623__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11378_ _11542_/A _11536_/A _11378_/C _11378_/D vssd1 vssd1 vccd1 vccd1 _11379_/B
+ sky130_fd_sc_hd__nand4_1
X_14166_ _14485_/CLK hold494/X vssd1 vssd1 vccd1 vccd1 hold493/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10329_ _10328_/B _10328_/C _10328_/A vssd1 vssd1 vccd1 vccd1 _10329_/Y sky130_fd_sc_hd__o21ai_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13489_/A hold31/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__and2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14097_ _15229_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 _14097_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13048_ hold265/A hold531/A _14618_/Q _13987_/Q _13091_/S _13098_/S1 vssd1 vssd1
+ vccd1 vccd1 _13048_/X sky130_fd_sc_hd__mux4_1
XANTENNA__08055__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A1 _13680_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12161__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14999_ _15254_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 _14999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07540_ hold633/X _13711_/A1 _07544_/S vssd1 vssd1 vccd1 vccd1 hold634/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_80_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08132__A1 _08564_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07471_ hold257/X _07473_/B vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__and2_1
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11812__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ _11288_/A1 _09209_/Y _09116_/X vssd1 vssd1 vccd1 vccd1 _12276_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12216__B1 _06926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13413__C1 _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _09138_/Y _09139_/X _09008_/X _09010_/X vssd1 vssd1 vccd1 vccd1 _09142_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12767__A1 _12917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_95_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__S0 _12365_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ _09119_/A _08957_/B _08954_/X vssd1 vssd1 vccd1 vccd1 _09073_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07310__B _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12519__A1 _12669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08023_ _08095_/A _08022_/B _07964_/A vssd1 vssd1 vccd1 vccd1 _08024_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13739__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold700 hold700/A vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout4 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout4/X sky130_fd_sc_hd__buf_4
XANTENNA__12614__S1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold711 hold711/A vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold722 hold722/A vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07737__S _07742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold733 hold733/A vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 hold744/A vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold755 hold755/A vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_153_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold777 hold777/A vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold788 hold788/A vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__xor2_1
Xhold799 hold799/A vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08141__B _08776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2101 _14766_/Q vssd1 vssd1 vccd1 vccd1 hold2101/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2112 _13207_/X vssd1 vssd1 vccd1 vccd1 _15071_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08925_ _10183_/A _09714_/A _11561_/A _09864_/A vssd1 vssd1 vccd1 vccd1 _09039_/A
+ sky130_fd_sc_hd__nand4_2
Xhold2123 _14362_/Q vssd1 vssd1 vccd1 vccd1 hold2123/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09699__A1 _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2134 _07123_/X vssd1 vssd1 vccd1 vccd1 _13933_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__B2 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2145 _13837_/Q vssd1 vssd1 vccd1 vccd1 hold2145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1400 _11900_/X vssd1 vssd1 vccd1 vccd1 _14721_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout576_A _15422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1411 _14546_/Q vssd1 vssd1 vccd1 vccd1 hold1411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2156 _07712_/X vssd1 vssd1 vccd1 vccd1 _14331_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1422 _07056_/X vssd1 vssd1 vccd1 vccd1 _13872_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2167 _14938_/Q vssd1 vssd1 vccd1 vccd1 _13499_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _14253_/Q vssd1 vssd1 vccd1 vccd1 hold1433/X sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ _08856_/A _14436_/Q _08856_/C vssd1 vssd1 vccd1 vccd1 _09087_/C sky130_fd_sc_hd__and3_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_168_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2178 _11742_/X vssd1 vssd1 vccd1 vccd1 _14536_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1444 _07199_/X vssd1 vssd1 vccd1 vccd1 _14006_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08371__A1 _08873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2189 _14653_/Q vssd1 vssd1 vccd1 vccd1 hold2189/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1455 _14355_/Q vssd1 vssd1 vccd1 vccd1 hold1455/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ hold1079/X _13745_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 _07807_/X sky130_fd_sc_hd__mux2_1
Xhold1466 _07609_/X vssd1 vssd1 vccd1 vccd1 _14233_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1477 _14724_/Q vssd1 vssd1 vccd1 vccd1 hold1477/X sky130_fd_sc_hd__dlygate4sd3_1
X_08787_ _08785_/X _08787_/B vssd1 vssd1 vccd1 vccd1 _08788_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout743_A _14953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1488 _11754_/X vssd1 vssd1 vccd1 vccd1 _14548_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _14311_/Q vssd1 vssd1 vccd1 vccd1 hold1499/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ hold735/X _13744_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 hold736/A sky130_fd_sc_hd__mux2_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09403__D _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__S0 _06943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11007__B _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ hold425/X _13741_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 hold426/A sky130_fd_sc_hd__mux2_1
XFILLER_0_95_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11722__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ _09408_/A _09408_/B _09408_/C vssd1 vssd1 vccd1 vccd1 _09411_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10680_ _11566_/A _15221_/Q vssd1 vssd1 vccd1 vccd1 _10681_/C sky130_fd_sc_hd__and2_1
XFILLER_0_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ _08526_/B _09337_/Y _09338_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _09339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_106_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _12692_/A1 _12347_/X _12349_/X vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ hold213/A _14328_/Q hold353/A _13988_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _11301_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12281_ _13168_/A _13448_/B vssd1 vssd1 vccd1 vccd1 _14930_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_160_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10862__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11232_ _11340_/A _15225_/Q vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07647__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14020_ _15384_/CLK hold402/X vssd1 vssd1 vccd1 vccd1 hold401/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09428__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12930__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ _11447_/A _11162_/B _10976_/A vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _10114_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ _10872_/A _10872_/B _10876_/B vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12143__C1 _13486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _10044_/B _10044_/C _10044_/A vssd1 vssd1 vccd1 vccd1 _10046_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__07890__B _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ _15242_/CLK _14922_/D vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfxtp_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09163__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2690 _14833_/Q vssd1 vssd1 vccd1 vccd1 hold2690/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _15254_/CLK _14853_/D vssd1 vssd1 vccd1 vccd1 _14853_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _15394_/CLK _13804_/D vssd1 vssd1 vccd1 vccd1 _13804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14784_ _15264_/CLK _14784_/D vssd1 vssd1 vccd1 vccd1 _14784_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13643__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ _14105_/Q _14098_/Q _11996_/C _14103_/Q vssd1 vssd1 vccd1 vccd1 _11997_/D
+ sky130_fd_sc_hd__or4b_1
X_13735_ hold427/X _13735_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold428/A sky130_fd_sc_hd__mux2_1
XFILLER_0_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _10932_/Y _10937_/Y _10946_/X _11509_/A _11511_/C1 vssd1 vssd1 vccd1 vccd1
+ _10948_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_196_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09862__A1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__B2 _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13666_ hold845/X _13666_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold846/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10878_ _10878_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13097__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07411__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ _15405_/CLK hold610/X vssd1 vssd1 vccd1 vccd1 hold609/A sky130_fd_sc_hd__dfxtp_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12642_/A1 _12616_/X _12642_/B1 vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__a21o_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12029__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ _11478_/B _11650_/B _13596_/X _13459_/A vssd1 vssd1 vccd1 vccd1 _13597_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15336_ _15340_/CLK _15336_/D vssd1 vssd1 vccd1 vccd1 _15336_/Q sky130_fd_sc_hd__dfxtp_1
X_12548_ hold225/A _14307_/Q _14598_/Q _13967_/Q _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12548_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09090__A2 _09925_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15267_ _15364_/CLK _15267_/D vssd1 vssd1 vccd1 vccd1 _15267_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _08175_/Y _12325_/B _12478_/X vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_112_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14218_ _15056_/CLK _14218_/D vssd1 vssd1 vccd1 vccd1 _14218_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09917__A2 _13395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15198_ _15199_/CLK _15198_/D vssd1 vssd1 vccd1 vccd1 _15198_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12382__C1 _13455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ _15080_/CLK _14149_/D vssd1 vssd1 vccd1 vccd1 _14149_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08050__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 _08065_/A vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06971_ _14083_/Q _14085_/Q _14091_/Q _14084_/Q vssd1 vssd1 vccd1 vccd1 _06972_/D
+ sky130_fd_sc_hd__or4b_1
XANTENNA__09225__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13021__S1 _13099_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _08712_/B vssd1 vssd1 vccd1 vccd1 _08710_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11807__S _11812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ _09690_/A _09690_/B _09690_/C vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__nand3_2
X_08641_ _08536_/B _08538_/B _08536_/A vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08572_ _08776_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nand2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ hold899/X _13727_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 hold900/A sky130_fd_sc_hd__mux2_1
XFILLER_0_193_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08200__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13323__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ _07454_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _14084_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07385_ _15346_/Q _07401_/A _14063_/Q _12294_/A _07382_/X vssd1 vssd1 vccd1 vccd1
+ _07385_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09124_ _09724_/D _09124_/B vssd1 vssd1 vccd1 vccd1 _09125_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_115_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09055_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__and3_2
XFILLER_0_103_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12373__S _12665_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ _08892_/A _10507_/A _11550_/A _08677_/A vssd1 vssd1 vccd1 vccd1 _08007_/C
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__12599__S0 _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09248__A _10142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold530 hold530/A vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 hold541/A vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08267__S1 _07815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold552 hold552/A vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12912__A1 _12949_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 hold563/A vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 hold574/A vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold585 hold585/A vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 hold596/A vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07991__A _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09957_ _10351_/A _10338_/D _09822_/A _09819_/Y vssd1 vssd1 vccd1 vccd1 _10065_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout860_A _07473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__C1 _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11717__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _08908_/A _09026_/B _09708_/B _09858_/C vssd1 vssd1 vccd1 vccd1 _08909_/C
+ sky130_fd_sc_hd__nand4_2
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09888_/A _09888_/B _09888_/C vssd1 vssd1 vccd1 vccd1 _09888_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__12402__A _13027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _07708_/X vssd1 vssd1 vccd1 vccd1 _14328_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__B1 _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 _14741_/Q vssd1 vssd1 vccd1 vccd1 hold1241/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12771__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1252 _07668_/X vssd1 vssd1 vccd1 vccd1 _14289_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ _08953_/B _08836_/X _08725_/X _08727_/Y vssd1 vssd1 vccd1 vccd1 _08840_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1263 _14330_/Q vssd1 vssd1 vccd1 vccd1 hold1263/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1274 _07658_/X vssd1 vssd1 vccd1 vccd1 _14279_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1285 _14312_/Q vssd1 vssd1 vccd1 vccd1 hold1285/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 _07635_/X vssd1 vssd1 vccd1 vccd1 _14258_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ hold1193/X _13737_/A1 _11861_/S vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12428__B1 _12953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__A1 _10741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ _10801_/A _10801_/B _10801_/C vssd1 vssd1 vccd1 vccd1 _10802_/B sky130_fd_sc_hd__and3_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12523__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ hold1397/X _13668_/A1 _11795_/S vssd1 vssd1 vccd1 vccd1 _11781_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13520_ _13668_/A1 hold1509/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09430__B _11586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _10733_/A _10733_/B vssd1 vssd1 vccd1 vccd1 _10734_/A sky130_fd_sc_hd__or2_1
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07231__A _15201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13451_ _09927_/B _13468_/A _13450_/Y _13409_/A vssd1 vssd1 vccd1 vccd1 _15219_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_211_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10663_ _10664_/A _10664_/B _10664_/C vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__and3_1
XFILLER_0_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07607__A0 _13746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ _13027_/A _12402_/B _12402_/C vssd1 vssd1 vccd1 vccd1 _12402_/X sky130_fd_sc_hd__and3_1
X_13382_ _13386_/A _13382_/B vssd1 vssd1 vccd1 vccd1 _15173_/D sky130_fd_sc_hd__and2_1
X_10594_ _11499_/B1 _10587_/Y _10589_/Y _10591_/Y _10593_/Y vssd1 vssd1 vccd1 vccd1
+ _10594_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15121_ _15127_/CLK _15121_/D vssd1 vssd1 vccd1 vccd1 _15121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12333_ _07912_/X _08636_/A _13140_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12334_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15052_ _15373_/CLK _15052_/D vssd1 vssd1 vccd1 vccd1 _15052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12264_ _13373_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _14913_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _15369_/CLK _14003_/D vssd1 vssd1 vccd1 vccd1 _14003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11215_ _11370_/A _11214_/B _11200_/Y vssd1 vssd1 vccd1 vccd1 _11215_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__12903__B2 _13195_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ _12128_/A _12195_/A2 _12194_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12195_/X
+ sky130_fd_sc_hd__o211a_1
X_11146_ _11146_/A _11146_/B _11146_/C vssd1 vssd1 vccd1 vccd1 _11148_/C sky130_fd_sc_hd__and3_1
XFILLER_0_208_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11077_ _11076_/B _11076_/C _11076_/A vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12667__B1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput150 in2[29] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__clkbuf_2
Xinput161 rst vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10028_ _10026_/X _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__and2b_1
X_14905_ _14992_/CLK _14905_/D vssd1 vssd1 vccd1 vccd1 _14905_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14836_ _14842_/CLK _14836_/D vssd1 vssd1 vccd1 vccd1 _14836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13616__C1 _07474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12514__S0 _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08099__B1 _10397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13092__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ _15377_/CLK hold864/X vssd1 vssd1 vccd1 vccd1 hold863/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11979_ hold1307/X _13668_/A1 _11993_/S vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10767__A _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13143__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__A1 _07879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ hold1497/X _13718_/A1 _13732_/S vssd1 vssd1 vccd1 vccd1 _13718_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ _15438_/CLK _14698_/D vssd1 vssd1 vccd1 vccd1 _14698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07941__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13649_ _07448_/A _13625_/C _13648_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15357_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07170_ _13671_/A1 hold2225/X _07181_/S vssd1 vssd1 vccd1 vccd1 _07170_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11598__A _11598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _15460_/CLK _15319_/D vssd1 vssd1 vccd1 vccd1 _15319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_120_clk clkbuf_4_8__f_clk/X vssd1 vssd1 vccd1 vccd1 _15188_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08403__C _08809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09811_ _09808_/Y _09964_/A _11335_/A _10166_/C vssd1 vssd1 vccd1 vccd1 _09964_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _09745_/C vssd1 vssd1 vccd1 vccd1 _09742_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06954_ _14029_/Q _14030_/Q vssd1 vssd1 vccd1 vccd1 _06962_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07316__A _15225_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _09673_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10133__A1 _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_187_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15072_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10133__B2 _11569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08491_/A _08492_/B _08621_/Y _08622_/X vssd1 vssd1 vccd1 vccd1 _08624_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11881__A1 _13735_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07750__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08760_/A _08555_/B vssd1 vssd1 vccd1 vccd1 _08555_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout441_A _08441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout539_A _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07506_ hold1625/X _13745_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 _07506_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07837__B1 _06959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ _08581_/A _08485_/C _08476_/Y vssd1 vssd1 vccd1 vccd1 _08487_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07932__S0 _08548_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10827__D _10827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07437_ _07437_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _14067_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12808__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ _15348_/Q _14061_/Q vssd1 vssd1 vccd1 vccd1 _07368_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12594__C1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ _09514_/A _09107_/B vssd1 vssd1 vccd1 vccd1 _09107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07299_ _07297_/Y _07299_/B vssd1 vssd1 vccd1 vccd1 _07320_/D sky130_fd_sc_hd__nand2b_1
XANTENNA__11492__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clkbuf_4_10__f_clk/X vssd1 vssd1 vccd1 vccd1 _15093_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07197__S _07198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ _08900_/A _08899_/B _08897_/X vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_142_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12116__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 hold360/A vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 hold371/A vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold382 hold382/A vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _11614_/A _11378_/D _11542_/B _11586_/A vssd1 vssd1 vccd1 vccd1 _11000_/X
+ sky130_fd_sc_hd__a22o_1
Xhold393 hold393/A vssd1 vssd1 vccd1 vccd1 hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__B2 _08760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout840 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _13041_/S sky130_fd_sc_hd__buf_6
Xfanout851 _13622_/C1 vssd1 vssd1 vccd1 vccd1 _13797_/C1 sky130_fd_sc_hd__buf_4
Xfanout862 _06946_/Y vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__buf_4
XFILLER_0_102_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout873 _13499_/A vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__buf_4
XANTENNA__12132__A _14877_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout884 _13390_/A vssd1 vssd1 vccd1 vccd1 _13389_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13310__A1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12113__A2 _12129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07226__A _15202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _12951_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _12952_/C sky130_fd_sc_hd__or2_1
XANTENNA__10124__A1 _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_178_clk clkbuf_leaf_0_clk/A vssd1 vssd1 vccd1 vccd1 _15042_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 _11847_/X vssd1 vssd1 vccd1 vccd1 _14670_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 _14316_/Q vssd1 vssd1 vccd1 vccd1 hold1071/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13662__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _13657_/A1 hold1993/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11902_/X sky130_fd_sc_hd__mux2_1
Xhold1082 _07632_/X vssd1 vssd1 vccd1 vccd1 _14255_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _13107_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _14963_/D sky130_fd_sc_hd__nor2_1
XANTENNA_200 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1093 _14113_/Q vssd1 vssd1 vccd1 vccd1 hold1093/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07660__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_222 _13375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _15261_/CLK hold856/X vssd1 vssd1 vccd1 vccd1 hold855/A sky130_fd_sc_hd__dfxtp_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ hold957/X hold2376/X _11845_/S vssd1 vssd1 vccd1 vccd1 hold958/A sky130_fd_sc_hd__mux2_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14552_ _14776_/CLK hold870/X vssd1 vssd1 vccd1 vccd1 hold869/A sky130_fd_sc_hd__dfxtp_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ hold1891/X _13651_/A1 _11779_/S vssd1 vssd1 vccd1 vccd1 _11764_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08057__A _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13651_/A1 hold2161/X _13518_/S vssd1 vssd1 vccd1 vccd1 _13503_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_138_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10715_ _10498_/X _10502_/C _10713_/Y _10714_/X vssd1 vssd1 vccd1 vccd1 _10717_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _14483_/CLK _14483_/D vssd1 vssd1 vccd1 vccd1 _14483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11695_ _14088_/Q _11729_/B _14090_/Q vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__or3_4
XANTENNA__11910__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13434_ _13440_/S _13434_/B vssd1 vssd1 vccd1 vccd1 _13434_/Y sky130_fd_sc_hd__nand2_1
X_10646_ _11564_/A _11623_/A _10646_/C _10646_/D vssd1 vssd1 vccd1 vccd1 _10646_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_183_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11388__B1 _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output193_A _15174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _13369_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _15156_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_102_clk clkbuf_leaf_88_clk/A vssd1 vssd1 vccd1 vccd1 _15242_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10577_ hold241/A hold961/A _14615_/Q _13984_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _10577_/X sky130_fd_sc_hd__mux4_1
X_15104_ _15116_/CLK _15104_/D vssd1 vssd1 vccd1 vccd1 _15104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _12316_/A vssd1 vssd1 vccd1 vccd1 _12316_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _13317_/A _13296_/B vssd1 vssd1 vccd1 vccd1 _15118_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15035_ _15457_/CLK _15035_/D vssd1 vssd1 vccd1 vccd1 _15035_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12741__S _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12247_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12983__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _14900_/Q _12178_/B vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__or2_1
XFILLER_0_208_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13138__A _13499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _11493_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13301__A1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_169_clk clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _15184_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12977__A _13102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14819_ _14840_/CLK _14819_/D vssd1 vssd1 vccd1 vccd1 _14819_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09808__A1 _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08340_ _08340_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08340_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11615__A1 _11567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ _14789_/Q hold709/A hold375/A _14725_/Q _07822_/S _12244_/S1 vssd1 vssd1
+ vccd1 vccd1 _08272_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12916__S _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07222_ _08677_/A _10873_/A vssd1 vssd1 vccd1 vccd1 _12254_/A sky130_fd_sc_hd__and2_1
XFILLER_0_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2740_A _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07153_ _13654_/A1 hold1525/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07084_ _13687_/A1 hold2187/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07084_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__C1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13747__S _13748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09526__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10354__A1 _11541_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_A _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ _08197_/A _07983_/X _07985_/X vssd1 vssd1 vccd1 vccd1 _07986_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_199_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09725_ _10033_/A _09726_/B _09726_/C _09726_/D vssd1 vssd1 vccd1 vccd1 _09727_/A
+ sky130_fd_sc_hd__a22oi_1
X_06937_ _06937_/A vssd1 vssd1 vccd1 vccd1 _06937_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10106__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _09533_/A _09532_/B _09532_/A vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10657__A2 _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07480__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ _08607_/A _08607_/B vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__xnor2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13056__B1 _08637_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09587_ _09587_/A _09587_/B vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__xnor2_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout823_A _12641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _13352_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12803__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08469_ _09008_/A _09860_/A vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _10323_/X _10328_/B _10498_/X _10499_/Y vssd1 vssd1 vccd1 vccd1 _10502_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11480_ _11111_/A _11111_/B _11290_/Y _11112_/A vssd1 vssd1 vccd1 vccd1 _11482_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ _11510_/A1 _10424_/Y _10426_/Y _10428_/Y _10430_/Y vssd1 vssd1 vccd1 vccd1
+ _10431_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_66_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _13150_/A _13150_/B vssd1 vssd1 vccd1 vccd1 _15015_/D sky130_fd_sc_hd__nor2_1
X_10362_ _10362_/A _10362_/B _10362_/C vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__nand3_2
XANTENNA__10593__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ hold2437/X _12129_/A2 _12100_/X _12037_/A vssd1 vssd1 vccd1 vccd1 _12101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13657__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ _10293_/A _10293_/B _10294_/B vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__and3_1
XFILLER_0_27_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ _13081_/A1 _13170_/B _08637_/Y vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07655__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ hold2471/X hold2550/X _12062_/S vssd1 vssd1 vccd1 vccd1 _12032_/X sky130_fd_sc_hd__mux2_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07882__C _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07210__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout670 hold2749/X vssd1 vssd1 vccd1 vccd1 _13708_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout681 hold103/X vssd1 vssd1 vccd1 vccd1 _13703_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout692 _15050_/Q vssd1 vssd1 vccd1 vccd1 _13730_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13983_ _15382_/CLK _13983_/D vssd1 vssd1 vccd1 vccd1 _13983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11905__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__A1 _13732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ hold437/A _13919_/Q _12941_/S vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ hold501/A _14128_/Q _12866_/S vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__mux2_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11206__A _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14604_ _15371_/CLK _14604_/D vssd1 vssd1 vccd1 vccd1 _14604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ hold1557/X _13703_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10110__A _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12796_ hold695/A _15280_/Q _15088_/Q _14381_/Q _12791_/S _12899_/S1 vssd1 vssd1
+ vccd1 vccd1 _12796_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_83_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _15400_/CLK _14535_/D vssd1 vssd1 vccd1 vccd1 _14535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11747_ _13700_/A1 hold1923/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__mux2_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14466_ _15437_/CLK _14466_/D vssd1 vssd1 vccd1 vccd1 _14466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _13742_/A1 hold1595/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11678_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13417_ hold443/X _13466_/A _13416_/Y _13178_/A vssd1 vssd1 vccd1 vccd1 hold444/A
+ sky130_fd_sc_hd__o211a_1
X_10629_ _10629_/A _10795_/B _10629_/C vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ _14397_/CLK hold382/X vssd1 vssd1 vccd1 vccd1 hold381/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08777__A1 _14950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ _13360_/A _13348_/B vssd1 vssd1 vccd1 vccd1 _15139_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10584__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08872__S1 _11306_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13279_ input132/X fanout6/X fanout4/X input100/X vssd1 vssd1 vccd1 vccd1 _13279_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10780__A _11580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08888__C _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ _15179_/CLK _15018_/D vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08250__A _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2508 hold2857/X vssd1 vssd1 vccd1 vccd1 _06905_/A sky130_fd_sc_hd__clkbuf_2
Xhold2519 _12125_/X vssd1 vssd1 vccd1 vccd1 _14874_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_166_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07840_ hold277/A _14034_/Q _14035_/Q vssd1 vssd1 vccd1 vccd1 _07841_/C sky130_fd_sc_hd__or3_1
XFILLER_0_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1807 _13923_/Q vssd1 vssd1 vccd1 vccd1 hold1807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1818 _07077_/X vssd1 vssd1 vccd1 vccd1 _13893_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__S0 _12741_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1829 _14374_/Q vssd1 vssd1 vccd1 vccd1 hold1829/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07771_ _11921_/A0 hold1977/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07771_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11815__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _09941_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08701__A1 _10033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__B2 _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _09439_/X _09441_/B vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15233__D _15233_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__B _11351_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _09514_/A _09372_/B vssd1 vssd1 vccd1 vccd1 _09372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_192_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ _08322_/B _08322_/C _08322_/A vssd1 vssd1 vccd1 vccd1 _08324_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_129_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08560__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08254_ _08252_/Y _08254_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07205_ hold675/X _13673_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold676/A sky130_fd_sc_hd__mux2_1
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ _14430_/Q _08441_/B vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__or2_1
XFILLER_0_132_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout404_A _11643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__A1 _08981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ _13737_/A1 hold1815/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07136_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10575__A1 _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__S1 _08868_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _13738_/A1 hold1381/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07067_/X sky130_fd_sc_hd__mux2_1
Xoutput240 _14444_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[20] sky130_fd_sc_hd__buf_12
Xoutput251 _14454_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[30] sky130_fd_sc_hd__buf_12
XFILLER_0_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput262 _14888_/Q vssd1 vssd1 vccd1 vccd1 out0[11] sky130_fd_sc_hd__buf_12
XFILLER_0_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput273 _14898_/Q vssd1 vssd1 vccd1 vccd1 out0[21] sky130_fd_sc_hd__buf_12
Xoutput284 _14908_/Q vssd1 vssd1 vccd1 vccd1 out0[31] sky130_fd_sc_hd__buf_12
XANTENNA_fanout773_A _11333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput295 _14857_/Q vssd1 vssd1 vccd1 vccd1 out1[12] sky130_fd_sc_hd__buf_12
XFILLER_0_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07969_ _07900_/B _13377_/B hold2377/X vssd1 vssd1 vccd1 vccd1 _07969_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11725__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _10126_/A _09708_/B _10126_/B _09858_/C vssd1 vssd1 vccd1 vccd1 _09709_/D
+ sky130_fd_sc_hd__nand4_4
X_10980_ _11563_/A _11569_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__and3_1
XFILLER_0_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09639_ _10244_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _09639_/X sky130_fd_sc_hd__or2_1
XFILLER_0_69_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07223__B _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ _12646_/X _12647_/X _12649_/X _12648_/X _12700_/S0 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12651_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_195_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ _11601_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11602_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12788__C1 _12988_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _08535_/A _08636_/A _13150_/B _13081_/A1 vssd1 vssd1 vccd1 vccd1 _12582_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08551__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14320_ _15380_/CLK hold560/X vssd1 vssd1 vccd1 vccd1 hold559/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _11532_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08208__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14251_ _15375_/CLK _14251_/D vssd1 vssd1 vccd1 vccd1 _14251_/Q sky130_fd_sc_hd__dfxtp_1
X_11463_ _11463_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11465_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08759__A1 _08989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13202_ _13404_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _15067_/D sky130_fd_sc_hd__and2_1
XANTENNA__13752__A1 _15459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ hold163/A hold627/A hold485/A _13983_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _10414_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09956__B1 _11514_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ _15184_/CLK hold130/X vssd1 vssd1 vccd1 vccd1 _14182_/Q sky130_fd_sc_hd__dfxtp_1
X_11394_ _11394_/A _11626_/A _11394_/C vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _13495_/A hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__and2_1
X_10345_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ hold1429/X hold823/X hold357/X hold1393/X _13066_/S _13068_/A1 vssd1 vssd1
+ vccd1 vccd1 _13064_/X sky130_fd_sc_hd__mux4_1
X_10276_ _11596_/A _11569_/B _14963_/Q _11577_/A vssd1 vssd1 vccd1 vccd1 _10277_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08070__A _12252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _12059_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _14820_/D sky130_fd_sc_hd__and2_1
XANTENNA__10105__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08220__D _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11818__A1 _15058_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13416__A _13466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13966_ _15077_/CLK _13966_/D vssd1 vssd1 vccd1 vccd1 _13966_/Q sky130_fd_sc_hd__dfxtp_1
X_12917_ _12917_/A1 _12916_/X _12917_/B1 vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_198_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13897_ _15434_/CLK _13897_/D vssd1 vssd1 vccd1 vccd1 _13897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12848_ hold201/A _14319_/Q _14610_/Q _13979_/Q _12915_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12848_/X sky130_fd_sc_hd__mux4_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12466__S _12466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ _13392_/B _13104_/A2 _12778_/X vssd1 vssd1 vccd1 vccd1 _12779_/X sky130_fd_sc_hd__a21o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08998__A1 _09846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10254__B1 _10255_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14518_ _15242_/CLK hold432/X vssd1 vssd1 vccd1 vccd1 hold431/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08998__B2 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ _15315_/CLK _14449_/D vssd1 vssd1 vccd1 vccd1 _14449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10006__B1 _10115_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 hold904/A vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 hold915/A vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10101__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 hold926/A vssd1 vssd1 vccd1 vccd1 hold926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 hold937/A vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold948 hold948/A vssd1 vssd1 vccd1 vccd1 hold948/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09990_ _09986_/X _09988_/Y _09831_/B _09833_/B vssd1 vssd1 vccd1 vccd1 _09990_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold959 hold959/A vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _08940_/B _08940_/C _08940_/A vssd1 vssd1 vccd1 vccd1 _08941_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2305 _14034_/Q vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold2316 _15328_/Q vssd1 vssd1 vccd1 vccd1 _07424_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold2703_A _15183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _14344_/Q _14248_/Q _14408_/Q _14120_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _08873_/B sky130_fd_sc_hd__mux4_1
Xhold2327 _13571_/X vssd1 vssd1 vccd1 vccd1 _15311_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2338 hold2862/X vssd1 vssd1 vccd1 vccd1 _07908_/A sky130_fd_sc_hd__buf_1
Xhold2349 _15034_/Q vssd1 vssd1 vccd1 vccd1 _07574_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 _11896_/X vssd1 vssd1 vccd1 vccd1 _14717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 _13989_/Q vssd1 vssd1 vccd1 vccd1 hold1615/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1626 _07506_/X vssd1 vssd1 vccd1 vccd1 _14134_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07823_ _12244_/S1 _07822_/X _08873_/A vssd1 vssd1 vccd1 vccd1 _07823_/X sky130_fd_sc_hd__a21o_1
Xhold1637 _14204_/Q vssd1 vssd1 vccd1 vccd1 hold1637/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1648 _07184_/X vssd1 vssd1 vccd1 vccd1 _13991_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1659 _15417_/Q vssd1 vssd1 vccd1 vccd1 hold1659/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13326__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09523__B _11536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _13659_/A1 hold457/X _07761_/S vssd1 vssd1 vccd1 vccd1 hold458/A sky130_fd_sc_hd__mux2_1
XFILLER_0_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07685_ hold345/X _13691_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold346/A sky130_fd_sc_hd__mux2_1
XFILLER_0_189_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_91_clk clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 _15258_/CLK sky130_fd_sc_hd__clkbuf_16
X_09424_ _09421_/A _09422_/X _09314_/B _09314_/Y vssd1 vssd1 vccd1 vccd1 _09461_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08438__B1 _09494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12234__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ _11104_/A _12277_/B _09354_/X vssd1 vssd1 vccd1 vccd1 _09355_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__07978__B _14426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A _08880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout619_A _15205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _08306_/A _08306_/B _08306_/C vssd1 vssd1 vccd1 vccd1 _08310_/A sky130_fd_sc_hd__nand3_1
X_09286_ _09285_/B _09285_/C _09285_/A vssd1 vssd1 vccd1 vccd1 _09288_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07110__A0 _15066_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08155__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10796__A1 _11563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10796__B2 _11594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ _08326_/B _08237_/B vssd1 vssd1 vccd1 vccd1 _08239_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08305__D _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ _08164_/Y _08165_/X _08166_/Y _08167_/Y _10397_/A vssd1 vssd1 vccd1 vccd1
+ _08174_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09402__A2 _11407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07119_ _13687_/A1 hold2005/X _07131_/S vssd1 vssd1 vccd1 vccd1 _07119_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08099_ _08097_/X _08098_/Y _10397_/A vssd1 vssd1 vccd1 vccd1 _08099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09961__A2_N _10338_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10130_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_63_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12124__B _12126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _10058_/Y _10059_/X _09841_/X _09896_/A vssd1 vssd1 vccd1 vccd1 _10061_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12396__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2850 _15357_/Q vssd1 vssd1 vccd1 vccd1 hold2850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2861 _15345_/Q vssd1 vssd1 vccd1 vccd1 hold2861/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13820_ _15191_/CLK _13820_/D vssd1 vssd1 vccd1 vccd1 _13820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__A _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13751_ hold2365/X _07812_/A _07391_/Y _13749_/Y _13750_/Y vssd1 vssd1 vccd1 vccd1
+ _13751_/X sky130_fd_sc_hd__a2111o_1
X_10963_ _11577_/A _14967_/Q vssd1 vssd1 vccd1 vccd1 _10964_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13670__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_clk _14581_/CLK vssd1 vssd1 vccd1 vccd1 _14419_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ _13102_/A _12702_/B _12702_/C vssd1 vssd1 vccd1 vccd1 _12702_/X sky130_fd_sc_hd__and3_1
XFILLER_0_74_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13682_ hold367/X _13715_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__mux2_1
X_10894_ _10893_/B _10893_/C _10893_/A vssd1 vssd1 vccd1 vccd1 _10894_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_167_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15421_ _15421_/CLK _15421_/D vssd1 vssd1 vccd1 vccd1 _15421_/Q sky130_fd_sc_hd__dfxtp_1
X_12633_ _15403_/Q _14538_/Q _14698_/Q _14762_/Q _12591_/S _12699_/S1 vssd1 vssd1
+ vccd1 vccd1 _12633_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12225__A1 _07900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12225__B2 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15352_ _15356_/CLK _15352_/D vssd1 vssd1 vccd1 vccd1 _15352_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12320__S1 _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ hold821/X hold1049/X hold899/X hold1223/X _12566_/S _12368_/A vssd1 vssd1
+ vccd1 vccd1 _12564_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_170_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08065__A _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ _15042_/CLK _14303_/D vssd1 vssd1 vccd1 vccd1 _14303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11515_ _07264_/A _11324_/X _07287_/Y vssd1 vssd1 vccd1 vccd1 _11515_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15283_ _15441_/CLK hold952/X vssd1 vssd1 vccd1 vccd1 hold951/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12495_ _12495_/A _12495_/B _12676_/A vssd1 vssd1 vccd1 vccd1 _12502_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12528__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234_ _15427_/CLK _14234_/D vssd1 vssd1 vccd1 vccd1 _14234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11446_ _11445_/A _11445_/B _11445_/C _11445_/D vssd1 vssd1 vccd1 vccd1 _11447_/C
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_145_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _14483_/CLK hold634/X vssd1 vssd1 vccd1 vccd1 hold633/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11377_ _11536_/A _11378_/C _11378_/D _11542_/A vssd1 vssd1 vccd1 vccd1 _11379_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13492_/A hold21/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__and2_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10328_ _10328_/A _10328_/B _10328_/C vssd1 vssd1 vccd1 vccd1 _10328_/X sky130_fd_sc_hd__or3_4
XANTENNA__07409__A _13501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _15229_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 _14096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ hold287/A hold413/A hold727/A _14746_/Q _13041_/S _13099_/S1 vssd1 vssd1
+ vccd1 vccd1 _13047_/X sky130_fd_sc_hd__mux4_1
X_10259_ _13708_/A1 _11514_/A2 _11514_/B1 _13196_/B _10257_/Y vssd1 vssd1 vccd1 vccd1
+ _10259_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13146__A _13381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ _15254_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 _14998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13949_ _15452_/CLK _13949_/D vssd1 vssd1 vccd1 vccd1 _13949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_clk clkbuf_leaf_76_clk/A vssd1 vssd1 vccd1 vccd1 _15289_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10475__B1 _11536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__S0 _08763_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ hold321/X _07475_/B vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07891__A1 _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12216__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__B1 _10107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09140_ _09008_/X _09010_/X _09138_/Y _09139_/X vssd1 vssd1 vccd1 vccd1 _09140_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12311__S1 _12365_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__A1 _13711_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__B2 _13199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2653_A _14979_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09071_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_154_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _08095_/A _08022_/B _07964_/A vssd1 vssd1 vccd1 vccd1 _08022_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_86_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08703__A _08926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 hold701/A vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold712 hold712/A vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout5 fanout6/A vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__buf_4
Xhold723 hold723/A vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold734 hold734/A vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 hold745/A vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold756 hold756/A vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 hold767/A vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap486 _07854_/Y vssd1 vssd1 vccd1 vccd1 _11474_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold778 hold778/A vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _10351_/A _11586_/B _09974_/A vssd1 vssd1 vccd1 vccd1 _09973_/Y sky130_fd_sc_hd__nand3_2
Xhold789 hold789/A vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10950__B2 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ _09714_/A _11561_/A _09864_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08926_/C
+ sky130_fd_sc_hd__a22o_1
Xhold2102 _11946_/X vssd1 vssd1 vccd1 vccd1 _14766_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2113 _14231_/Q vssd1 vssd1 vccd1 vccd1 hold2113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2124 _07746_/X vssd1 vssd1 vccd1 vccd1 _14362_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09699__A2 _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2135 _13922_/Q vssd1 vssd1 vccd1 vccd1 hold2135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07753__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1401 _14591_/Q vssd1 vssd1 vccd1 vccd1 hold1401/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2146 _07020_/X vssd1 vssd1 vccd1 vccd1 _13837_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1412 _11752_/X vssd1 vssd1 vccd1 vccd1 _14546_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ _14436_/Q _08856_/C _08856_/A vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__a21oi_1
Xhold2157 _15412_/Q vssd1 vssd1 vccd1 vccd1 hold2157/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout471_A _12128_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1423 _14222_/Q vssd1 vssd1 vccd1 vccd1 hold1423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2168 _13499_/X vssd1 vssd1 vccd1 vccd1 _15258_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold2179 _13874_/Q vssd1 vssd1 vccd1 vccd1 hold2179/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _07630_/X vssd1 vssd1 vccd1 vccd1 _14253_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1445 _14755_/Q vssd1 vssd1 vccd1 vccd1 hold1445/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A _10425_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1456 _07736_/X vssd1 vssd1 vccd1 vccd1 _14355_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07806_ hold309/X _13744_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 hold310/A sky130_fd_sc_hd__mux2_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08786_ _08785_/B _08785_/C _08785_/A vssd1 vssd1 vccd1 vccd1 _08787_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1467 _14217_/Q vssd1 vssd1 vccd1 vccd1 hold1467/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1478 _11903_/X vssd1 vssd1 vccd1 vccd1 _14724_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 _13867_/Q vssd1 vssd1 vccd1 vccd1 hold1489/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_211_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12455__A1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ hold2143/X _13743_/A1 _07742_/S vssd1 vssd1 vccd1 vccd1 _07737_/X sky130_fd_sc_hd__mux2_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_A _11390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_clk clkbuf_leaf_92_clk/A vssd1 vssd1 vccd1 vccd1 _14866_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07989__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__S1 _12700_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11007__C _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ hold1251/X _13740_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 _07668_/X sky130_fd_sc_hd__mux2_1
X_09407_ _09539_/B _09406_/C _09406_/A vssd1 vssd1 vccd1 vccd1 _09408_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_137_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12207__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07599_ _13705_/A1 hold1703/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07599_/X sky130_fd_sc_hd__mux2_1
X_09338_ _09338_/A _12256_/A vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ _09269_/A _09269_/B vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12834__S _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ _13594_/A _13591_/A2 _11289_/Y _11299_/Y _13459_/A vssd1 vssd1 vccd1 vccd1
+ _11300_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09709__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _13168_/A _13446_/B vssd1 vssd1 vccd1 vccd1 _14929_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__B _15222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ _11231_/A _11231_/B vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09428__B _09708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07229__A _11606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _11447_/A _11162_/B _10976_/A vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__nor3b_2
XANTENNA__09139__A1 _09138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13665__S _13666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _10280_/B _10111_/X _10000_/X _10003_/B vssd1 vssd1 vccd1 vccd1 _10114_/B
+ sky130_fd_sc_hd__a211oi_2
X_11093_ _11093_/A _11093_/B vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07663__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A _10002_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _10044_/A _10044_/B _10044_/C vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__and3_2
X_14921_ _15242_/CLK _14921_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12694__A1 _12700_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2680 _14442_/Q vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09163__B _09979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2691 _15050_/Q vssd1 vssd1 vccd1 vccd1 hold2691/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _15254_/CLK _14852_/D vssd1 vssd1 vccd1 vccd1 _14852_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13803_ _14754_/CLK _13803_/D vssd1 vssd1 vccd1 vccd1 _13803_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1990 _11732_/X vssd1 vssd1 vccd1 vccd1 _14526_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14783_ _14783_/CLK _14783_/D vssd1 vssd1 vccd1 vccd1 _14783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11995_ _14099_/Q _11995_/B vssd1 vssd1 vccd1 vccd1 _11997_/C sky130_fd_sc_hd__or2_1
XFILLER_0_97_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15354_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10457__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ hold723/X _13734_/A1 _13748_/S vssd1 vssd1 vccd1 vccd1 hold724/A sky130_fd_sc_hd__mux2_1
X_10946_ _11510_/A1 _10939_/Y _10941_/Y _10943_/Y _10945_/Y vssd1 vssd1 vccd1 vccd1
+ _10946_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07873__A1 _15342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13665_ hold581/X _13665_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold582/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ _10651_/A _10650_/B _10648_/X vssd1 vssd1 vccd1 vccd1 _10887_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12616_ _14342_/Q _14246_/Q _12735_/S vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__mux2_1
X_15404_ _15441_/CLK hold910/X vssd1 vssd1 vccd1 vccd1 hold909/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07411__B _07411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _14454_/Q _13636_/B vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__or2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15335_ _15354_/CLK _15335_/D vssd1 vssd1 vccd1 vccd1 _15335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ hold665/A _14502_/Q hold569/A _14726_/Q _12441_/S _12674_/S1 vssd1 vssd1
+ vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_108_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15432_/CLK _15266_/D vssd1 vssd1 vccd1 vccd1 _15266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ _13690_/A1 _12329_/B _12953_/B1 _13178_/B vssd1 vssd1 vccd1 vccd1 _12478_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_3 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14217_ _15405_/CLK _14217_/D vssd1 vssd1 vccd1 vccd1 _14217_/Q sky130_fd_sc_hd__dfxtp_1
X_11429_ _11578_/A _14970_/Q vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_112_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09338__B _12256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15197_ _15424_/CLK _15197_/D vssd1 vssd1 vccd1 vccd1 _15197_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _15437_/CLK hold900/X vssd1 vssd1 vccd1 vccd1 hold899/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10932__A1 _11493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06970_ _06972_/C _06970_/B vssd1 vssd1 vccd1 vccd1 _11997_/B sky130_fd_sc_hd__or2_1
X_14079_ _14083_/CLK hold128/X vssd1 vssd1 vccd1 vccd1 _14079_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09225__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__A2 _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08984__S0 _09239_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ _08640_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08642_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ _08571_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__or2_1
XANTENNA__12437__A1 _12674_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_clk clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 _15425_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09302__A1 _10185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11823__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07522_ hold1929/X _13693_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07522_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2770_A _14492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07453_ _07453_/A _13317_/A vssd1 vssd1 vccd1 vccd1 _14083_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07384_ _15347_/Q _07402_/A _14061_/Q _07439_/A _07383_/X vssd1 vssd1 vccd1 vccd1
+ _07387_/C sky130_fd_sc_hd__o221a_1
XFILLER_0_162_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09123_ _09846_/B _09724_/C _09724_/D _11580_/A vssd1 vssd1 vccd1 vccd1 _09125_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10963__A _11577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07748__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _09051_/Y _09052_/X _08933_/Y _08935_/X vssd1 vssd1 vccd1 vccd1 _09055_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08005_ _08677_/A _08892_/A _10507_/A _11550_/A vssd1 vssd1 vccd1 vccd1 _08007_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_170_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09248__B _10142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12599__S1 _12599_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 hold520/A vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold531 hold531/A vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold542 hold542/A vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold553 hold553/A vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold564 hold564/A vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 hold575/A vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold586 hold586/A vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold597/A vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ _13673_/A1 _11514_/A2 _11514_/B1 _13194_/B _09954_/Y vssd1 vssd1 vccd1 vccd1
+ _09956_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_60_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07483__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ _09026_/B _09708_/B _09858_/C _08908_/A vssd1 vssd1 vccd1 vccd1 _08909_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09264__A _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09888_/A _09888_/B _09888_/C vssd1 vssd1 vccd1 vccd1 _09887_/X sky130_fd_sc_hd__and3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout853_A _13622_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 _07709_/X vssd1 vssd1 vccd1 vccd1 _14329_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A1 _09979_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 _14804_/Q vssd1 vssd1 vccd1 vccd1 hold1231/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__B2 _10183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _08725_/X _08727_/Y _08953_/B _08836_/X vssd1 vssd1 vccd1 vccd1 _08838_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08975__S0 _08990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1242 _11920_/X vssd1 vssd1 vccd1 vccd1 _14741_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1253 _14687_/Q vssd1 vssd1 vccd1 vccd1 hold1253/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12771__S1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1264 _07711_/X vssd1 vssd1 vccd1 vccd1 _14330_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1275 _15391_/Q vssd1 vssd1 vccd1 vccd1 hold1275/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _07692_/X vssd1 vssd1 vccd1 vccd1 _14312_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _08992_/A1 _08762_/Y _08764_/Y _08766_/Y _08768_/Y vssd1 vssd1 vccd1 vccd1
+ _08769_/X sky130_fd_sc_hd__o32a_1
Xhold1297 _14763_/Q vssd1 vssd1 vccd1 vccd1 hold1297/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12428__B2 _13176_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _14955_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11733__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ _10801_/A _10801_/B _10801_/C vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__a21oi_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12523__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12979__A2 _13104_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ hold585/X _13519_/A0 _11795_/S vssd1 vssd1 vccd1 vccd1 hold586/A sky130_fd_sc_hd__mux2_1
XFILLER_0_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ _10558_/A _10558_/B _10557_/A vssd1 vssd1 vccd1 vccd1 _10733_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09430__C _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07231__B _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13450_ _13450_/A _13450_/B vssd1 vssd1 vccd1 vccd1 _13450_/Y sky130_fd_sc_hd__nand2_1
X_10662_ _10491_/A _10491_/C _10491_/B vssd1 vssd1 vccd1 vccd1 _10664_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _12676_/A _12401_/B vssd1 vssd1 vccd1 vccd1 _12402_/C sky130_fd_sc_hd__or2_1
XFILLER_0_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ _13381_/A _13381_/B vssd1 vssd1 vccd1 vccd1 _15172_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_180_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10873__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _11507_/A _10592_/X _11499_/B1 vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15120_ _15127_/CLK _15120_/D vssd1 vssd1 vccd1 vccd1 _15120_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07658__S _07660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12332_ _13374_/B _12330_/B _12327_/Y _12331_/Y _12328_/X vssd1 vssd1 vccd1 vccd1
+ _13140_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15441_/CLK _15051_/D vssd1 vssd1 vccd1 vccd1 _15051_/Q sky130_fd_sc_hd__dfxtp_1
X_12263_ _13381_/A _13412_/B vssd1 vssd1 vccd1 vccd1 _14912_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11167__A1 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ _14569_/CLK hold304/X vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__dfxtp_1
X_11214_ _11370_/A _11214_/B _11200_/Y vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__nor3b_2
XANTENNA__13561__C1 _13565_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12903__A2 _13103_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ _14908_/Q _12194_/B vssd1 vssd1 vccd1 vccd1 _12194_/X sky130_fd_sc_hd__or2_1
XANTENNA__11908__S _11911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _11146_/A _11146_/B _11146_/C vssd1 vssd1 vccd1 vccd1 _11148_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11076_ _11076_/A _11076_/B _11076_/C vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__or3_1
XANTENNA__12667__A1 _12692_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12211__S0 _12198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_clk_A clkbuf_leaf_99_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput140 in2[1] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07421__A_N _07812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput151 in2[2] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_2
X_10027_ _10024_/X _10025_/Y _09863_/X _09865_/X vssd1 vssd1 vccd1 vccd1 _10028_/B
+ sky130_fd_sc_hd__a211o_1
X_14904_ _14992_/CLK _14904_/D vssd1 vssd1 vccd1 vccd1 _14904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07406__B _13317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _14842_/CLK _14835_/D vssd1 vssd1 vccd1 vccd1 _14835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12419__A1 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_clk clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 _14783_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12514__S1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13092__A1 _13092_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ hold1581/X _13519_/A0 _11993_/S vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__mux2_1
X_14766_ _15439_/CLK _14766_/D vssd1 vssd1 vccd1 vccd1 _14766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13143__B _13143_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_152_clk_A clkbuf_4_3__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ hold1661/X _12329_/A _13732_/S vssd1 vssd1 vccd1 vccd1 _13717_/X sky130_fd_sc_hd__mux2_1
X_10929_ hold259/A hold317/A hold703/A _13986_/Q _10930_/S0 _10930_/S1 vssd1 vssd1
+ vccd1 vccd1 _10929_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11642__A2 _11641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14697_ _15440_/CLK _14697_/D vssd1 vssd1 vccd1 vccd1 _14697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07941__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ input57/X _13648_/B vssd1 vssd1 vccd1 vccd1 _13648_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_32_clk_A clkbuf_4_6__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ _09919_/B _13586_/B _13578_/X _13579_/C1 vssd1 vssd1 vccd1 vccd1 _13579_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_167_clk_A clkbuf_4_2__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__B _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ _15423_/CLK _15318_/D vssd1 vssd1 vccd1 vccd1 _15318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08253__A _08253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_clk_A clkbuf_4_5__f_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _15250_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12450__S0 _12644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ _09661_/A _10166_/C _09808_/Y _09964_/A vssd1 vssd1 vccd1 vccd1 _09812_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11818__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09741_ _09741_/A _09741_/B _09599_/B vssd1 vssd1 vccd1 vccd1 _09745_/C sky130_fd_sc_hd__nor3b_2
X_06953_ _06953_/A _14028_/Q _14029_/Q _06952_/X vssd1 vssd1 vccd1 vccd1 _06953_/X
+ sky130_fd_sc_hd__or4bb_1
XANTENNA__12202__S0 _12237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15236__D _15236_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_105_clk_A _14581_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ _09578_/A _09577_/B _09575_/X vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07316__B _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08623_ _08491_/A _08492_/B _08621_/Y _08622_/X vssd1 vssd1 vccd1 vccd1 _08623_/Y
+ sky130_fd_sc_hd__a211oi_2
Xclkbuf_leaf_19_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15226_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08989_/A _08551_/X _08553_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08555_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07505_ hold759/X _13744_/A1 _07509_/S vssd1 vssd1 vccd1 vccd1 hold760/A sky130_fd_sc_hd__mux2_1
X_08485_ _08476_/Y _08581_/A _08485_/C vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12830__A1 _13080_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout434_A _07778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _08964_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _14066_/D sky130_fd_sc_hd__and2_1
XANTENNA__07932__S1 _08548_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10693__A _10873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A _09860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ _15348_/Q _14061_/Q vssd1 vssd1 vccd1 vccd1 _07367_/X sky130_fd_sc_hd__or2_1
XANTENNA__12384__S _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _14282_/Q _14218_/Q _14154_/Q _14472_/Q _09239_/S0 _09239_/S1 vssd1 vssd1
+ vccd1 vccd1 _09107_/B sky130_fd_sc_hd__mux4_1
XANTENNA__07478__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07298_ _11620_/B _11594_/B vssd1 vssd1 vccd1 vccd1 _07299_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11492__S1 _11501_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _09037_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold350 hold350/A vssd1 vssd1 vccd1 vccd1 hold350/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 hold361/A vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/A vssd1 vssd1 vccd1 vccd1 hold383/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__S _11728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 hold394/A vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout830 _12791_/S vssd1 vssd1 vccd1 vccd1 _12741_/S sky130_fd_sc_hd__buf_8
Xfanout841 _12964_/S0 vssd1 vssd1 vccd1 vccd1 _13091_/S sky130_fd_sc_hd__buf_4
Xfanout852 _13622_/C1 vssd1 vssd1 vccd1 vccd1 _13409_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09939_ hold551/A hold951/A hold837/A _14384_/Q _11306_/S0 _11306_/S1 vssd1 vssd1
+ vccd1 vccd1 _09939_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_205_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout863 _13397_/A vssd1 vssd1 vccd1 vccd1 _13396_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout874 _13501_/A vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__buf_2
Xfanout885 _13107_/A vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__buf_4
XANTENNA__07226__B _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _12946_/X _12947_/X _12949_/X _12948_/X _12950_/S0 _13100_/S1 vssd1 vssd1
+ vccd1 vccd1 _12951_/B sky130_fd_sc_hd__mux4_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10124__A2 _11594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _07588_/X vssd1 vssd1 vccd1 vccd1 _14212_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 _14251_/Q vssd1 vssd1 vccd1 vccd1 hold1061/X sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _13656_/A1 hold1353/X _11911_/S vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__mux2_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1072 _07696_/X vssd1 vssd1 vccd1 vccd1 _14316_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 _14122_/Q vssd1 vssd1 vccd1 vccd1 hold1083/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _13106_/A1 _13162_/B _13031_/B1 vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__o21a_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _07485_/X vssd1 vssd1 vccd1 vccd1 _14113_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12559__S _12566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _15192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _15292_/CLK hold558/X vssd1 vssd1 vccd1 vccd1 hold557/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_223 _13375_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ hold453/X _13719_/A1 _11845_/S vssd1 vssd1 vccd1 vccd1 hold454/A sky130_fd_sc_hd__mux2_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08338__A _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07242__A _10356_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09373__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _15416_/CLK hold828/X vssd1 vssd1 vccd1 vccd1 hold827/A sky130_fd_sc_hd__dfxtp_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _13716_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10713_/B _10713_/C _10713_/A vssd1 vssd1 vccd1 vccd1 _10714_/X sky130_fd_sc_hd__o21a_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13502_/A _13502_/B vssd1 vssd1 vccd1 vccd1 _13502_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__08772__S _10949_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14775_/CLK _14482_/D vssd1 vssd1 vccd1 vccd1 _14482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ _06903_/A _13792_/A2 _11693_/X _07475_/B vssd1 vssd1 vccd1 vccd1 _14492_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13433_ _13541_/A _13433_/B vssd1 vssd1 vccd1 vccd1 _15210_/D sky130_fd_sc_hd__and2_1
XFILLER_0_180_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10645_ _11564_/A _11623_/A _10646_/C _10646_/D vssd1 vssd1 vccd1 vccd1 _10645_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_153_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11388__A1 _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11388__B2 _11588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13364_ _13369_/A _13364_/B vssd1 vssd1 vccd1 vccd1 _15155_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08073__A _08312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10576_ _06914_/A _13586_/B _10575_/Y _13409_/A vssd1 vssd1 vccd1 vccd1 _10576_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_output186_A _15196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ _15116_/CLK _15103_/D vssd1 vssd1 vccd1 vccd1 _15103_/Q sky130_fd_sc_hd__dfxtp_1
X_12315_ _12311_/X _12312_/X _12314_/X _12313_/X _12366_/A _06944_/A vssd1 vssd1 vccd1
+ vccd1 _12316_/A sky130_fd_sc_hd__mux4_1
X_13295_ input73/X fanout2/X _13294_/X vssd1 vssd1 vccd1 vccd1 _13296_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10108__A _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15034_ _15289_/CLK _15034_/D vssd1 vssd1 vccd1 vccd1 _15034_/Q sky130_fd_sc_hd__dfxtp_1
X_12246_ hold853/A _13927_/Q _15428_/Q _13895_/Q _12237_/S _12231_/A vssd1 vssd1 vccd1
+ vccd1 _12247_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12888__A1 _12917_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ hold2553/X _12195_/A2 _12176_/X _13491_/A vssd1 vssd1 vccd1 vccd1 _12177_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12983__S1 _13024_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__A1 _14947_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ hold629/A hold797/A hold489/A _14135_/Q _11506_/S0 _11506_/S1 vssd1 vssd1
+ vccd1 vccd1 _11129_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_78_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _11351_/B _11614_/B _11586_/B _11541_/A vssd1 vssd1 vccd1 vccd1 _11062_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13154__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818_ _14844_/CLK _14818_/D vssd1 vssd1 vccd1 vccd1 _14818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12499__S0 _12460_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__A2 _09809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08248__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07819__A1 _12243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__A2 _15227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12812__A1 _06942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14749_ _15426_/CLK _14749_/D vssd1 vssd1 vccd1 vccd1 _14749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08270_ _15366_/Q _15269_/Q hold527/A hold457/A _07816_/S _07815_/A vssd1 vssd1 vccd1
+ vccd1 _08270_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07332_/B sky130_fd_sc_hd__inv_2
XANTENNA_hold2566_A _15355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__A _13389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ _13653_/A1 hold1547/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07152_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12671__S0 _12735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07083_ _13719_/A1 hold2115/X _07096_/S vssd1 vssd1 vccd1 vccd1 _07083_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _15313_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12423__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__A1 _13396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13329__A _13338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11000__B1 _11542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B _10338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12233__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__S1 _13074_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__A2 _11561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07985_ _08201_/A _07984_/X _12201_/C1 vssd1 vssd1 vccd1 vccd1 _07985_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout384_A _11895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _10115_/A _10115_/B _09724_/C _09724_/D vssd1 vssd1 vccd1 vccd1 _09726_/D
+ sky130_fd_sc_hd__nand4_1
X_06936_ hold277/X vssd1 vssd1 vccd1 vccd1 hold278/A sky130_fd_sc_hd__inv_2
XANTENNA__11303__A1 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _10351_/A _10166_/C _09537_/A _09534_/X vssd1 vssd1 vccd1 vccd1 _09754_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout551_A _15423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__S _11283_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08606_ _08699_/B _08606_/B vssd1 vssd1 vccd1 vccd1 _08607_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout649_A _15198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09586_ _09587_/A _09587_/B vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__and2_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13056__A1 _07355_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ _08437_/A _08434_/Y _08436_/B vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12803__B2 _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout816_A _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07997__A _08065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _08468_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ hold17/X _07473_/B vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__and2_1
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08399_ _09164_/A _09712_/A _08468_/A _08400_/D vssd1 vssd1 vccd1 vccd1 _08411_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12567__B1 _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _10244_/A _10429_/X _10430_/B1 vssd1 vssd1 vccd1 vccd1 _10430_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07001__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _10524_/B _10360_/C _10360_/A vssd1 vssd1 vccd1 vccd1 _10362_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12100_ _14990_/Q _12126_/B _12126_/C _12128_/D vssd1 vssd1 vccd1 vccd1 _12100_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13080_ _13080_/A1 _13079_/X hold2771/X vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__a21oi_1
X_10292_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10294_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12414__S0 _12459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12031_ _12037_/A _12031_/B vssd1 vssd1 vccd1 vccd1 _14828_/D sky130_fd_sc_hd__and2_1
XANTENNA__13239__A _15353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout660 _15065_/Q vssd1 vssd1 vccd1 vccd1 _13745_/A1 sky130_fd_sc_hd__buf_4
Xfanout671 _13740_/A1 vssd1 vssd1 vccd1 vccd1 _13674_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13673__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout682 _13735_/A1 vssd1 vssd1 vccd1 vccd1 _13669_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13295__A1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout693 _15050_/Q vssd1 vssd1 vccd1 vccd1 _13664_/A1 sky130_fd_sc_hd__clkbuf_4
X_13982_ _15090_/CLK _13982_/D vssd1 vssd1 vccd1 vccd1 _13982_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09499__B1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07671__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ hold419/A hold983/A hold331/A _14774_/Q _12916_/S _12949_/S1 vssd1 vssd1
+ vccd1 vccd1 _12933_/X sky130_fd_sc_hd__mux4_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09171__B _09858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ hold593/A _14224_/Q hold691/A hold729/A _12866_/S _13074_/S1 vssd1 vssd1
+ vccd1 vccd1 _12864_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14603_ _15367_/CLK _14603_/D vssd1 vssd1 vccd1 vccd1 _14603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11206__B _11623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ hold1257/X _13669_/A1 _11828_/S vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__mux2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12795_ _12795_/A _12795_/B _12951_/A vssd1 vssd1 vccd1 vccd1 _12802_/B sky130_fd_sc_hd__or3b_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10110__B _14961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11921__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ _13732_/A1 hold1573/X _11761_/S vssd1 vssd1 vccd1 vccd1 _11746_/X sky130_fd_sc_hd__mux2_1
X_14534_ _15045_/CLK hold750/X vssd1 vssd1 vccd1 vccd1 hold749/A sky130_fd_sc_hd__dfxtp_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _13708_/A1 hold1927/X _11684_/S vssd1 vssd1 vccd1 vccd1 _11677_/X sky130_fd_sc_hd__mux2_1
X_14465_ _15360_/CLK _14465_/D vssd1 vssd1 vccd1 vccd1 _14465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10628_ _10795_/A _10627_/C _10627_/A vssd1 vssd1 vccd1 vccd1 _10629_/C sky130_fd_sc_hd__a21o_1
X_13416_ _13466_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_181_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14396_ _15392_/CLK _14396_/D vssd1 vssd1 vccd1 vccd1 _14396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13347_ _13360_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _15138_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10559_ _10560_/A _10560_/B _10560_/C vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07985__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13278_ _13287_/A _13278_/B vssd1 vssd1 vccd1 vccd1 _15112_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10780__B _11578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ _15179_/CLK _15017_/D vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13149__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _12243_/A _12229_/B vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_209_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09346__B _09346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08250__B _08250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2509 _14988_/Q vssd1 vssd1 vccd1 vccd1 hold2509/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_166_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1808 _07110_/X vssd1 vssd1 vccd1 vccd1 _13923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1819 _14246_/Q vssd1 vssd1 vccd1 vccd1 hold1819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12708__S1 _12749_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07770_ _13675_/A1 hold1975/X _07777_/S vssd1 vssd1 vccd1 vccd1 _07770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07581__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12494__C1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08701__A2 _08809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _09437_/Y _09438_/X _09252_/X _09254_/X vssd1 vssd1 vccd1 vccd1 _09441_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13038__A1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09371_ _14671_/Q _13944_/Q hold427/A _13912_/Q _10429_/S0 _10429_/S1 vssd1 vssd1
+ vccd1 vccd1 _09372_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13589__A2 _13591_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11831__S _11845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _08322_/A _08322_/B _08322_/C vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold2850_A _15357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08254_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08560__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07204_ hold621/X _13705_/A1 _07214_/S vssd1 vssd1 vccd1 vccd1 hold622/A sky130_fd_sc_hd__mux2_1
XFILLER_0_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08184_ _09494_/A1 _08114_/Y _08183_/X vssd1 vssd1 vccd1 vccd1 _08184_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07135_ _13736_/A1 hold2083/X _07147_/S vssd1 vssd1 vccd1 vccd1 _07135_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10575__A2 _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__S _07761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07066_ _13671_/A1 hold1387/X _07077_/S vssd1 vssd1 vccd1 vccd1 _07066_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput230 _14435_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[11] sky130_fd_sc_hd__buf_12
Xoutput241 _14445_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[21] sky130_fd_sc_hd__buf_12
XANTENNA_fanout599_A _09676_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput252 _14455_/Q vssd1 vssd1 vccd1 vccd1 imemreq_addr[31] sky130_fd_sc_hd__buf_12
Xoutput263 _14889_/Q vssd1 vssd1 vccd1 vccd1 out0[12] sky130_fd_sc_hd__buf_12
Xoutput274 _14899_/Q vssd1 vssd1 vccd1 vccd1 out0[22] sky130_fd_sc_hd__buf_12
XANTENNA__12947__S1 _13098_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput285 _14880_/Q vssd1 vssd1 vccd1 vccd1 out0[3] sky130_fd_sc_hd__buf_12
XFILLER_0_11_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput296 _14858_/Q vssd1 vssd1 vccd1 vccd1 out1[13] sky130_fd_sc_hd__buf_12
XFILLER_0_96_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07968_ _07951_/Y _07967_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _13377_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07491__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09707_ _09708_/B _10126_/B _09858_/C _10126_/A vssd1 vssd1 vccd1 vccd1 _09709_/C
+ sky130_fd_sc_hd__a22o_1
X_06919_ _06919_/A vssd1 vssd1 vccd1 vccd1 _07402_/A sky130_fd_sc_hd__inv_2
X_07899_ _07899_/A _07899_/B vssd1 vssd1 vccd1 vccd1 _07899_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__11307__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09638_ _14801_/Q _14513_/Q hold615/A _14737_/Q _09795_/S0 _09795_/S1 vssd1 vssd1
+ vccd1 vccd1 _09639_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13029__A1 _11102_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09569_ _09714_/A _09714_/C _09864_/D _09571_/A vssd1 vssd1 vccd1 vccd1 _09573_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _11600_/A _11600_/B vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09102__C1 _10430_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ _12327_/A _12579_/X _12577_/X vssd1 vssd1 vccd1 vccd1 _13150_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12883__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ _11340_/A _15227_/Q _11366_/X _11368_/Y vssd1 vssd1 vccd1 vccd1 _11532_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08551__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11042__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _15374_/CLK hold546/X vssd1 vssd1 vccd1 vccd1 hold545/A sky130_fd_sc_hd__dfxtp_1
X_11462_ _11463_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11462_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ _13404_/A _13201_/B vssd1 vssd1 vccd1 vccd1 _15066_/D sky130_fd_sc_hd__and2_1
XANTENNA__13668__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _13584_/A _13797_/A2 _10412_/X _13797_/C1 vssd1 vssd1 vccd1 vccd1 _10413_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ _15184_/CLK hold136/X vssd1 vssd1 vccd1 vccd1 _14181_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09500__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10881__A _11517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11393_ _11392_/B _11392_/C _11392_/A vssd1 vssd1 vccd1 vccd1 _11394_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09956__B2 _13194_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _13495_/A hold153/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__and2_1
XANTENNA__07666__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13063_ _06943_/A _13058_/X _13062_/X _14491_/Q vssd1 vssd1 vccd1 vccd1 _13070_/A
+ sky130_fd_sc_hd__o211a_1
X_10275_ _11577_/A _11596_/A _11569_/B _11563_/B vssd1 vssd1 vccd1 vccd1 _10275_/X
+ sky130_fd_sc_hd__and4_1
X_12014_ hold2634/X hold2659/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11916__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12601__A _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout490 _12128_/B vssd1 vssd1 vccd1 vccd1 _12126_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13416__B _13416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ _15264_/CLK _13965_/D vssd1 vssd1 vccd1 vccd1 _13965_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ _14354_/Q _14258_/Q _12916_/S vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__mux2_1
X_13896_ _15429_/CLK _13896_/D vssd1 vssd1 vccd1 vccd1 _13896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ _14802_/Q _14514_/Q hold323/A hold865/A _12841_/S _06942_/A vssd1 vssd1 vccd1
+ vccd1 _12847_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13440__A1 _12277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12778_ _13735_/A1 _13103_/A2 _13078_/B1 _13190_/B vssd1 vssd1 vccd1 vccd1 _12778_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12874__S0 _12866_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__A1 _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__A2 _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__B _13151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517_ _15382_/CLK _14517_/D vssd1 vssd1 vccd1 vccd1 _14517_/Q sky130_fd_sc_hd__dfxtp_1
X_11729_ _14088_/Q _11729_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__or3_4
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ _15423_/CLK _14448_/D vssd1 vssd1 vccd1 vccd1 _14448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10006__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10006__B2 _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__B1 _11623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14379_ _15375_/CLK _14379_/D vssd1 vssd1 vccd1 vccd1 _14379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold905 hold905/A vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 hold916/A vssd1 vssd1 vccd1 vccd1 hold916/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10101__S1 _10930_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold927 hold927/A vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 hold938/A vssd1 vssd1 vccd1 vccd1 hold938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 hold949/A vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08940_ _08940_/A _08940_/B _08940_/C vssd1 vssd1 vccd1 vccd1 _08940_/Y sky130_fd_sc_hd__nand3_2
XANTENNA_hold2529_A _14069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12703__B1 _13078_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2306 _06937_/Y vssd1 vssd1 vccd1 vccd1 _07459_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_209_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2317 _14027_/Q vssd1 vssd1 vccd1 vccd1 _07452_/A sky130_fd_sc_hd__dlygate4sd3_1
X_08871_ _15426_/Q _08871_/B vssd1 vssd1 vccd1 vccd1 _08871_/Y sky130_fd_sc_hd__nor2_1
Xhold2328 _15163_/Q vssd1 vssd1 vccd1 vccd1 hold2328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2339 _13539_/X vssd1 vssd1 vccd1 vccd1 _15295_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1605 _14792_/Q vssd1 vssd1 vccd1 vccd1 hold1605/X sky130_fd_sc_hd__dlygate4sd3_1
X_07822_ hold763/A _14719_/Q _07822_/S vssd1 vssd1 vccd1 vccd1 _07822_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11826__S _11828_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1616 _07181_/X vssd1 vssd1 vccd1 vccd1 _13989_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13259__A1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1627 _13975_/Q vssd1 vssd1 vccd1 vccd1 hold1627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1638 _07580_/X vssd1 vssd1 vccd1 vccd1 _14204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 _14319_/Q vssd1 vssd1 vccd1 vccd1 hold1649/X sky130_fd_sc_hd__dlygate4sd3_1
X_07753_ _13724_/A1 hold1985/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07753_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_211_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11127__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ hold333/X _13657_/A1 _07693_/S vssd1 vssd1 vccd1 vccd1 hold334/A sky130_fd_sc_hd__mux2_1
XFILLER_0_189_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09423_ _09314_/B _09314_/Y _09421_/A _09422_/X vssd1 vssd1 vccd1 vccd1 _09461_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09354_ _08256_/A _13359_/B _09352_/X _09353_/Y vssd1 vssd1 vccd1 vccd1 _09354_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09635__B1 _11303_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08305_ _10507_/A _08776_/B _09026_/B _09138_/A vssd1 vssd1 vccd1 vccd1 _08306_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__10245__A1 _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09285_ _09285_/A _09285_/B _09285_/C vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08155__B _08702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout514_A _10252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10796__A2 _11606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__A1 _13715_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ _08093_/A _08158_/X _08289_/A vssd1 vssd1 vccd1 vccd1 _08237_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09938__A1 _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ _08164_/Y _08165_/X _08166_/Y vssd1 vssd1 vccd1 vccd1 _08167_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__S _07493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__B1 _06943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ _13719_/A1 hold975/X _07131_/S vssd1 vssd1 vccd1 vccd1 hold976/A sky130_fd_sc_hd__mux2_1
X_08098_ _07965_/Y _08024_/B _08022_/Y vssd1 vssd1 vccd1 vccd1 _08098_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout883_A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07049_ _13654_/A1 hold2175/X _07061_/S vssd1 vssd1 vccd1 vccd1 _07049_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ _09841_/X _09896_/A _10058_/Y _10059_/X vssd1 vssd1 vccd1 vccd1 _10060_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09797__S0 _10429_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__S _11745_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2840 _15336_/Q vssd1 vssd1 vccd1 vccd1 hold2840/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09714__B _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2851 _15303_/Q vssd1 vssd1 vccd1 vccd1 hold2851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2862 _15295_/Q vssd1 vssd1 vccd1 vccd1 hold2862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__B _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _14969_/Q _10781_/B _10961_/X vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__a21bo_1
X_13750_ _13750_/A _13750_/B vssd1 vssd1 vccd1 vccd1 _13750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12701_ _12951_/A _12701_/B vssd1 vssd1 vccd1 vccd1 _12702_/C sky130_fd_sc_hd__or2_1
XFILLER_0_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10893_ _10893_/A _10893_/B _10893_/C vssd1 vssd1 vccd1 vccd1 _11038_/B sky130_fd_sc_hd__or3_2
X_13681_ hold953/X _13681_/A1 _13682_/S vssd1 vssd1 vccd1 vccd1 hold954/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15420_ _15457_/CLK hold784/X vssd1 vssd1 vccd1 vccd1 hold783/A sky130_fd_sc_hd__dfxtp_1
X_12632_ _13150_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _14953_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_195_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07250__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__A1 _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15351_ _15351_/CLK _15351_/D vssd1 vssd1 vccd1 vccd1 _15351_/Q sky130_fd_sc_hd__dfxtp_1
X_12563_ _12366_/A _12558_/X _12562_/X _06944_/A vssd1 vssd1 vccd1 vccd1 _12570_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14302_ _15265_/CLK _14302_/D vssd1 vssd1 vccd1 vccd1 _14302_/Q sky130_fd_sc_hd__dfxtp_1
X_11514_ _13715_/A1 _11514_/A2 _11514_/B1 _13203_/B _11512_/Y vssd1 vssd1 vccd1 vccd1
+ _11514_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_163_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12494_ _12644_/A1 _12489_/X _12493_/X _12675_/S1 vssd1 vssd1 vccd1 vccd1 _12495_/B
+ sky130_fd_sc_hd__o211a_1
X_15282_ _15379_/CLK _15282_/D vssd1 vssd1 vccd1 vccd1 _15282_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12608__S0 _12441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11445_ _11445_/A _11445_/B _11445_/C _11445_/D vssd1 vssd1 vccd1 vccd1 _11593_/B
+ sky130_fd_sc_hd__or4_2
X_14233_ _15456_/CLK _14233_/D vssd1 vssd1 vccd1 vccd1 _14233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10095__S0 _10930_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _14775_/CLK _14164_/D vssd1 vssd1 vccd1 vccd1 _14164_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08601__A1 _09008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ _11376_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08601__B2 _09858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10327_ _10326_/B _10326_/C _10326_/A vssd1 vssd1 vccd1 vccd1 _10328_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13115_ _13489_/A hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__and2_1
X_14095_ _15229_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _14095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07409__B _07409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13033__S0 _13041_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _15387_/Q _15290_/Q hold753/A _14391_/Q _13091_/S _13098_/S1 vssd1 vssd1
+ vccd1 vccd1 _13046_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10258_ hold2737/X input17/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13196_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_56_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12161__A1 hold2562/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10189_ _10189_/A _10189_/B _10189_/C vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13146__B _13146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14997_ _15004_/CLK hold154/X vssd1 vssd1 vccd1 vccd1 _14997_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08117__B1 _12201_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08668__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13948_ _15062_/CLK _13948_/D vssd1 vssd1 vccd1 vccd1 _13948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10475__A1 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10475__B2 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__S1 _08763_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10786__A _11597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ _15375_/CLK _13879_/D vssd1 vssd1 vccd1 vccd1 _13879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13162__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07891__A2 _08075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__S0 _12841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__A _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10227__A1 _11288_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B1 _14969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__A2 _11514_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09070_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _08091_/B _08020_/B _08020_/C vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold2646_A _15166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08279__S0 _07816_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08703__B _09437_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 hold702/A vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/A vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10086__S0 _10087_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout6 fanout6/A vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__buf_4
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 hold724/A vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1__f_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold735 hold735/A vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 hold746/A vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 hold757/A vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold768 hold768/A vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _14941_/Q _11586_/B vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__nand2_1
Xhold779 hold779/A vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12940__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13024__S0 _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__A2 _12260_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08923_ _09435_/A _09860_/A _08775_/X _08776_/X _14950_/Q vssd1 vssd1 vccd1 vccd1
+ _08928_/A sky130_fd_sc_hd__a32o_1
Xhold2103 _13862_/Q vssd1 vssd1 vccd1 vccd1 hold2103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2114 _07607_/X vssd1 vssd1 vccd1 vccd1 _14231_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12688__C1 _06944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2125 _13943_/Q vssd1 vssd1 vccd1 vccd1 hold2125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold2136 _07109_/X vssd1 vssd1 vccd1 vccd1 _13922_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2147 _13900_/Q vssd1 vssd1 vccd1 vccd1 hold2147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1402 _11766_/X vssd1 vssd1 vccd1 vccd1 _14591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _14509_/Q vssd1 vssd1 vccd1 vccd1 hold1413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2158 _13706_/X vssd1 vssd1 vccd1 vccd1 _15412_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ _08854_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _13355_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12241__A _12241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1424 _07598_/X vssd1 vssd1 vccd1 vccd1 _14222_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08451__S0 _07822_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12481__A1_N _08179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2169 _15279_/Q vssd1 vssd1 vccd1 vccd1 hold2169/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 _14009_/Q vssd1 vssd1 vccd1 vccd1 hold1435/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1446 _11935_/X vssd1 vssd1 vccd1 vccd1 _14755_/D sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ hold2213/X _13743_/A1 _07810_/S vssd1 vssd1 vccd1 vccd1 _07805_/X sky130_fd_sc_hd__mux2_1
X_08785_ _08785_/A _08785_/B _08785_/C vssd1 vssd1 vccd1 vccd1 _08785_/X sky130_fd_sc_hd__and3_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1457 _14227_/Q vssd1 vssd1 vccd1 vccd1 hold1457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _07593_/X vssd1 vssd1 vccd1 vccd1 _14217_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout464_A _07045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1479 _13956_/Q vssd1 vssd1 vccd1 vccd1 hold1479/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ hold1455/X _11921_/A0 _07742_/S vssd1 vssd1 vccd1 vccd1 _07736_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13652__A1 _13652_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07667_ hold593/X _13739_/A1 _07676_/S vssd1 vssd1 vccd1 vccd1 hold594/A sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout631_A _15202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11007__D _11537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout729_A _14959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09406_ _09406_/A _09539_/B _09406_/C vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07598_ _13737_/A1 hold1423/X _07609_/S vssd1 vssd1 vccd1 vccd1 _07598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_165_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09337_ _09762_/C _09337_/B vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _09269_/B _09269_/A vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08219_ _09661_/A _09138_/A vssd1 vssd1 vccd1 vccd1 _08222_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ _09199_/A _09199_/B vssd1 vssd1 vccd1 vccd1 _09201_/B sky130_fd_sc_hd__or2_1
XANTENNA__09709__B _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11231_/A _11231_/B vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11320__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10926__C1 _07390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _11160_/B _11160_/C _11160_/A vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12470__C_N _12676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _10000_/X _10003_/B _10280_/B _10111_/X vssd1 vssd1 vccd1 vccd1 _10114_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_207_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11092_ _11093_/B _11093_/A vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12143__A1 hold2621/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _10042_/A _10042_/B _10042_/C vssd1 vssd1 vccd1 vccd1 _10044_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14920_ _15367_/CLK _14920_/D vssd1 vssd1 vccd1 vccd1 _14920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09444__B _10110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07245__A _09864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2670 _15142_/Q vssd1 vssd1 vccd1 vccd1 hold2670/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold2681 _09496_/X vssd1 vssd1 vccd1 vccd1 _14442_/D sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ _15254_/CLK _14851_/D vssd1 vssd1 vccd1 vccd1 _14851_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2692 _14434_/Q vssd1 vssd1 vccd1 vccd1 _08542_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13681__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13802_ _14595_/CLK hold930/X vssd1 vssd1 vccd1 vccd1 hold929/A sky130_fd_sc_hd__dfxtp_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1980 _07125_/X vssd1 vssd1 vccd1 vccd1 _13935_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13643__A1 _08345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1991 _14239_/Q vssd1 vssd1 vccd1 vccd1 hold1991/X sky130_fd_sc_hd__dlygate4sd3_1
X_14782_ _15427_/CLK _14782_/D vssd1 vssd1 vccd1 vccd1 _14782_/Q sky130_fd_sc_hd__dfxtp_1
X_11994_ _14100_/Q _14101_/Q _14102_/Q _14104_/Q vssd1 vssd1 vccd1 vccd1 _11995_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_187_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10457__A1 _11573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10457__B2 _11590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ hold395/X _15053_/Q _13748_/S vssd1 vssd1 vccd1 vccd1 hold396/A sky130_fd_sc_hd__mux2_1
X_10945_ _11493_/A _10944_/X _11510_/A1 vssd1 vssd1 vccd1 vccd1 _10945_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13664_ hold459/X _13664_/A1 _13666_/S vssd1 vssd1 vccd1 vccd1 hold460/A sky130_fd_sc_hd__mux2_1
X_10876_ _10876_/A _10876_/B vssd1 vssd1 vccd1 vccd1 _10893_/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ _15440_/CLK _15403_/D vssd1 vssd1 vccd1 vccd1 _15403_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11406__B1 _11570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12615_ hold1865/X hold1527/X _12641_/S vssd1 vssd1 vccd1 vccd1 _12615_/X sky130_fd_sc_hd__mux2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ _11291_/B _11650_/B _13594_/X _13459_/A vssd1 vssd1 vccd1 vccd1 _15323_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11501__S0 _11501_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15340_/CLK _15334_/D vssd1 vssd1 vccd1 vccd1 _15334_/Q sky130_fd_sc_hd__dfxtp_1
X_12546_ hold339/A _15270_/Q hold889/A _14371_/Q _12665_/S _12668_/A1 vssd1 vssd1
+ vccd1 vccd1 _12546_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_124_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ _15265_/CLK _15265_/D vssd1 vssd1 vccd1 vccd1 _15265_/Q sky130_fd_sc_hd__dfxtp_1
X_12477_ _13027_/A _12477_/B _12477_/C vssd1 vssd1 vccd1 vccd1 _12477_/X sky130_fd_sc_hd__and3_1
XANTENNA_4 _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__B1 _13031_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _15079_/CLK _14216_/D vssd1 vssd1 vccd1 vccd1 _14216_/Q sky130_fd_sc_hd__dfxtp_1
X_11428_ _11580_/A _14971_/Q vssd1 vssd1 vccd1 vccd1 _11430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _15196_/CLK _15196_/D vssd1 vssd1 vccd1 vccd1 _15196_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12382__A1 _07919_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__B2 _13081_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ _11518_/B _11358_/C _11358_/A vssd1 vssd1 vccd1 vccd1 _11359_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12760__S _12916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14147_ _15360_/CLK _14147_/D vssd1 vssd1 vccd1 vccd1 _14147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14078_ _15356_/CLK _14078_/D vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13157__A _13389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ _11102_/Y _13104_/A2 _13028_/X vssd1 vssd1 vccd1 vccd1 _13029_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12061__A _12063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_leaf_7_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__S1 _09239_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08570_ _08569_/B _08569_/C _08569_/A vssd1 vssd1 vccd1 vccd1 _08570_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07521_ hold1827/X _13725_/A1 _07528_/S vssd1 vssd1 vccd1 vccd1 _07521_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09370__A _10426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09302__A2 _09709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ _07452_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__and2_1
XANTENNA__12000__S _12062_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold2763_A _15186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07321__C _07321_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ _07437_/A _14059_/Q _07403_/A _15348_/Q vssd1 vssd1 vccd1 vccd1 _07383_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12935__S _12941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _09164_/A _09979_/C _09037_/A _09034_/X vssd1 vssd1 vccd1 vccd1 _09198_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10963__B _14967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _08933_/Y _08935_/X _09051_/Y _09052_/X vssd1 vssd1 vccd1 vccd1 _09055_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08004_ hold2372/X _12260_/A2 _12259_/A1 _13176_/B _08002_/Y vssd1 vssd1 vccd1 vccd1
+ _08004_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold510 hold510/A vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09248__C _10126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold521 hold521/A vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold532 hold532/A vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold543 hold543/A vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold554 hold554/A vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/A vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold576 hold576/A vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_204_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07764__S _07777_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 hold587/A vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 hold598/A vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ hold2727/X input15/X _10949_/S vssd1 vssd1 vccd1 vccd1 _13194_/B sky130_fd_sc_hd__mux2_2
XANTENNA_fanout581_A _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _09661_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__and2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09264__B _09726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _09886_/A _09886_/B _09886_/C vssd1 vssd1 vccd1 vccd1 _09888_/C sky130_fd_sc_hd__nand3_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _07749_/X vssd1 vssd1 vccd1 vccd1 _14365_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _15407_/Q vssd1 vssd1 vccd1 vccd1 hold1221/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A2 _15209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 _11985_/X vssd1 vssd1 vccd1 vccd1 _14804_/D sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ _08725_/X _08727_/Y _08953_/B _08836_/X vssd1 vssd1 vccd1 vccd1 _08840_/A
+ sky130_fd_sc_hd__a211oi_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08975__S1 _08990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1243 _14706_/Q vssd1 vssd1 vccd1 vccd1 hold1243/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout846_A _13477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1254 _11865_/X vssd1 vssd1 vccd1 vccd1 _14687_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1265 _14283_/Q vssd1 vssd1 vccd1 vccd1 hold1265/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1276 _13685_/X vssd1 vssd1 vccd1 vccd1 _15391_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1287 _13881_/Q vssd1 vssd1 vccd1 vccd1 hold1287/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08981_/A _08767_/X _08992_/A1 vssd1 vssd1 vccd1 vccd1 _08768_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12428__A2 _12329_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1298 _11943_/X vssd1 vssd1 vccd1 vccd1 _14763_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ hold461/X _13725_/A1 _07726_/S vssd1 vssd1 vccd1 vccd1 hold462/A sky130_fd_sc_hd__mux2_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08699_ _08699_/A _08699_/B vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11315__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10730_ _10730_/A _10730_/B vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07004__S _07010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10661_ _10660_/B _10660_/C _10660_/A vssd1 vssd1 vccd1 vccd1 _10664_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ _12396_/X _12397_/X _12399_/X _12398_/X _12644_/A1 _12675_/S1 vssd1 vssd1
+ vccd1 vccd1 _12401_/B sky130_fd_sc_hd__mux4_1
X_13380_ _13381_/A _13380_/B vssd1 vssd1 vccd1 vccd1 _15171_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10592_ hold819/A hold827/A _14711_/Q _14775_/Q _11316_/S0 _11316_/S1 vssd1 vssd1
+ vccd1 vccd1 _10592_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10873__B _15224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _13172_/B _12953_/B1 _12329_/X vssd1 vssd1 vccd1 vccd1 _12331_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15050_ _15179_/CLK _15050_/D vssd1 vssd1 vccd1 vccd1 _15050_/Q sky130_fd_sc_hd__dfxtp_1
X_12262_ _13481_/A _12262_/B vssd1 vssd1 vccd1 vccd1 _14911_/D sky130_fd_sc_hd__and2_1
XFILLER_0_160_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ _11212_/A _11212_/B _11212_/C vssd1 vssd1 vccd1 vccd1 _11214_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08568__B1 _12259_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14001_ _15080_/CLK hold892/X vssd1 vssd1 vccd1 vccd1 hold891/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13676__S _13682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__A2 _08526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ hold2610/X _12195_/A2 _12192_/X _13489_/A vssd1 vssd1 vccd1 vccd1 _12193_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08663__S0 _08868_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07674__S _07676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _11596_/A _14967_/Q vssd1 vssd1 vccd1 vccd1 _11146_/C sky130_fd_sc_hd__and2_1
XFILLER_0_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11075_ _11076_/A _11076_/B _11076_/C vssd1 vssd1 vccd1 vccd1 _11075_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__10127__B1 _10827_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput130 in2[10] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12211__S1 _12211_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput141 in2[20] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__clkbuf_2
Xinput152 in2[30] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__clkbuf_2
X_10026_ _09863_/X _09865_/X _10024_/X _10025_/Y vssd1 vssd1 vccd1 vccd1 _10026_/X
+ sky130_fd_sc_hd__o211a_1
X_14903_ _14987_/CLK _14903_/D vssd1 vssd1 vccd1 vccd1 _14903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output229_A _14434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__S _11927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _14842_/CLK _14834_/D vssd1 vssd1 vccd1 vccd1 _14834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13616__A1 _07431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13424__B _13424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _15056_/CLK _14765_/D vssd1 vssd1 vccd1 vccd1 _14765_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ hold937/X _13666_/A1 _11977_/S vssd1 vssd1 vccd1 vccd1 hold938/A sky130_fd_sc_hd__mux2_1
XFILLER_0_129_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11225__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13716_ _13716_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13716_/Y sky130_fd_sc_hd__nor2_4
X_10928_ _14451_/Q _13591_/A2 _10920_/Y hold2358/X _13409_/A vssd1 vssd1 vccd1 vccd1
+ _10928_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14696_ _15042_/CLK _14696_/D vssd1 vssd1 vccd1 vccd1 _14696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _08535_/A _13792_/A2 _13646_/X _07474_/B vssd1 vssd1 vccd1 vccd1 _15356_/D
+ sky130_fd_sc_hd__o211a_1
X_10859_ _11037_/B _10857_/X _10673_/A _10673_/Y vssd1 vssd1 vccd1 vccd1 _10900_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_128_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12052__A0 hold2535/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__A _08535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ _14445_/Q _13590_/B vssd1 vssd1 vccd1 vccd1 _13578_/X sky130_fd_sc_hd__or2_1
XFILLER_0_171_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ _15423_/CLK _15317_/D vssd1 vssd1 vccd1 vccd1 _15317_/Q sky130_fd_sc_hd__dfxtp_1
X_12529_ _13382_/B _12325_/B _12528_/X vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15248_ _15248_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__S _12491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15179_ _15179_/CLK _15179_/D vssd1 vssd1 vccd1 vccd1 _15179_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09220__A1 _09918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09220__B2 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12450__S1 _12675_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07584__S _07593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__C _10283_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A2 _13394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A1 _13687_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09739_/B _09739_/C _09739_/A vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__a21oi_1
X_06952_ _14027_/Q _14026_/Q _14030_/Q vssd1 vssd1 vccd1 vccd1 _06952_/X sky130_fd_sc_hd__and3_1
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10304__A _11605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
.ends


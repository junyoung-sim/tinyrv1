// This is the unpowered netlist.
module Proc (clk,
    dmemreq_type,
    dmemreq_val,
    imemreq_val,
    rst,
    dmemreq_addr,
    dmemreq_wdata,
    dmemresp_rdata,
    imemreq_addr,
    imemresp_data,
    in0,
    in1,
    in2,
    out0,
    out1,
    out2);
 input clk;
 output dmemreq_type;
 output dmemreq_val;
 output imemreq_val;
 input rst;
 output [31:0] dmemreq_addr;
 output [31:0] dmemreq_wdata;
 input [31:0] dmemresp_rdata;
 output [31:0] imemreq_addr;
 input [31:0] imemresp_data;
 input [31:0] in0;
 input [31:0] in1;
 input [31:0] in2;
 output [31:0] out0;
 output [31:0] out1;
 output [31:0] out2;

 wire net895;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire \ctrl.c2d_rf_waddr_W[0] ;
 wire \ctrl.c2d_rf_waddr_W[1] ;
 wire \ctrl.c2d_rf_waddr_W[2] ;
 wire \ctrl.c2d_rf_waddr_W[3] ;
 wire \ctrl.c2d_rf_waddr_W[4] ;
 wire \ctrl.d2c_inst[0] ;
 wire \ctrl.d2c_inst[10] ;
 wire \ctrl.d2c_inst[11] ;
 wire \ctrl.d2c_inst[12] ;
 wire \ctrl.d2c_inst[13] ;
 wire \ctrl.d2c_inst[14] ;
 wire \ctrl.d2c_inst[15] ;
 wire \ctrl.d2c_inst[16] ;
 wire \ctrl.d2c_inst[17] ;
 wire \ctrl.d2c_inst[18] ;
 wire \ctrl.d2c_inst[19] ;
 wire \ctrl.d2c_inst[1] ;
 wire \ctrl.d2c_inst[20] ;
 wire \ctrl.d2c_inst[21] ;
 wire \ctrl.d2c_inst[22] ;
 wire \ctrl.d2c_inst[23] ;
 wire \ctrl.d2c_inst[24] ;
 wire \ctrl.d2c_inst[25] ;
 wire \ctrl.d2c_inst[26] ;
 wire \ctrl.d2c_inst[27] ;
 wire \ctrl.d2c_inst[28] ;
 wire \ctrl.d2c_inst[29] ;
 wire \ctrl.d2c_inst[2] ;
 wire \ctrl.d2c_inst[30] ;
 wire \ctrl.d2c_inst[31] ;
 wire \ctrl.d2c_inst[3] ;
 wire \ctrl.d2c_inst[4] ;
 wire \ctrl.d2c_inst[5] ;
 wire \ctrl.d2c_inst[6] ;
 wire \ctrl.d2c_inst[7] ;
 wire \ctrl.d2c_inst[8] ;
 wire \ctrl.d2c_inst[9] ;
 wire \ctrl.inst_M[0] ;
 wire \ctrl.inst_M[10] ;
 wire \ctrl.inst_M[11] ;
 wire \ctrl.inst_M[12] ;
 wire \ctrl.inst_M[13] ;
 wire \ctrl.inst_M[14] ;
 wire \ctrl.inst_M[1] ;
 wire \ctrl.inst_M[20] ;
 wire \ctrl.inst_M[21] ;
 wire \ctrl.inst_M[22] ;
 wire \ctrl.inst_M[23] ;
 wire \ctrl.inst_M[24] ;
 wire \ctrl.inst_M[25] ;
 wire \ctrl.inst_M[26] ;
 wire \ctrl.inst_M[27] ;
 wire \ctrl.inst_M[28] ;
 wire \ctrl.inst_M[29] ;
 wire \ctrl.inst_M[2] ;
 wire \ctrl.inst_M[30] ;
 wire \ctrl.inst_M[31] ;
 wire \ctrl.inst_M[3] ;
 wire \ctrl.inst_M[4] ;
 wire \ctrl.inst_M[5] ;
 wire \ctrl.inst_M[6] ;
 wire \ctrl.inst_M[7] ;
 wire \ctrl.inst_M[8] ;
 wire \ctrl.inst_M[9] ;
 wire \ctrl.inst_W[0] ;
 wire \ctrl.inst_W[12] ;
 wire \ctrl.inst_W[13] ;
 wire \ctrl.inst_W[14] ;
 wire \ctrl.inst_W[1] ;
 wire \ctrl.inst_W[20] ;
 wire \ctrl.inst_W[21] ;
 wire \ctrl.inst_W[22] ;
 wire \ctrl.inst_W[23] ;
 wire \ctrl.inst_W[24] ;
 wire \ctrl.inst_W[25] ;
 wire \ctrl.inst_W[26] ;
 wire \ctrl.inst_W[27] ;
 wire \ctrl.inst_W[28] ;
 wire \ctrl.inst_W[29] ;
 wire \ctrl.inst_W[2] ;
 wire \ctrl.inst_W[30] ;
 wire \ctrl.inst_W[31] ;
 wire \ctrl.inst_W[3] ;
 wire \ctrl.inst_W[4] ;
 wire \ctrl.inst_W[5] ;
 wire \ctrl.inst_W[6] ;
 wire \ctrl.inst_X[0] ;
 wire \ctrl.inst_X[10] ;
 wire \ctrl.inst_X[11] ;
 wire \ctrl.inst_X[12] ;
 wire \ctrl.inst_X[13] ;
 wire \ctrl.inst_X[14] ;
 wire \ctrl.inst_X[1] ;
 wire \ctrl.inst_X[20] ;
 wire \ctrl.inst_X[21] ;
 wire \ctrl.inst_X[22] ;
 wire \ctrl.inst_X[23] ;
 wire \ctrl.inst_X[24] ;
 wire \ctrl.inst_X[25] ;
 wire \ctrl.inst_X[26] ;
 wire \ctrl.inst_X[27] ;
 wire \ctrl.inst_X[28] ;
 wire \ctrl.inst_X[29] ;
 wire \ctrl.inst_X[2] ;
 wire \ctrl.inst_X[30] ;
 wire \ctrl.inst_X[31] ;
 wire \ctrl.inst_X[3] ;
 wire \ctrl.inst_X[4] ;
 wire \ctrl.inst_X[5] ;
 wire \ctrl.inst_X[6] ;
 wire \ctrl.inst_X[7] ;
 wire \ctrl.inst_X[8] ;
 wire \ctrl.inst_X[9] ;
 wire \ctrl.val_D ;
 wire \ctrl.val_DX.q ;
 wire \ctrl.val_M ;
 wire \ctrl.val_MW.q ;
 wire \dpath.RF.R[0][0] ;
 wire \dpath.RF.R[0][10] ;
 wire \dpath.RF.R[0][11] ;
 wire \dpath.RF.R[0][12] ;
 wire \dpath.RF.R[0][13] ;
 wire \dpath.RF.R[0][14] ;
 wire \dpath.RF.R[0][15] ;
 wire \dpath.RF.R[0][16] ;
 wire \dpath.RF.R[0][17] ;
 wire \dpath.RF.R[0][18] ;
 wire \dpath.RF.R[0][19] ;
 wire \dpath.RF.R[0][1] ;
 wire \dpath.RF.R[0][20] ;
 wire \dpath.RF.R[0][21] ;
 wire \dpath.RF.R[0][22] ;
 wire \dpath.RF.R[0][23] ;
 wire \dpath.RF.R[0][24] ;
 wire \dpath.RF.R[0][25] ;
 wire \dpath.RF.R[0][26] ;
 wire \dpath.RF.R[0][27] ;
 wire \dpath.RF.R[0][28] ;
 wire \dpath.RF.R[0][29] ;
 wire \dpath.RF.R[0][2] ;
 wire \dpath.RF.R[0][30] ;
 wire \dpath.RF.R[0][31] ;
 wire \dpath.RF.R[0][3] ;
 wire \dpath.RF.R[0][4] ;
 wire \dpath.RF.R[0][5] ;
 wire \dpath.RF.R[0][6] ;
 wire \dpath.RF.R[0][7] ;
 wire \dpath.RF.R[0][8] ;
 wire \dpath.RF.R[0][9] ;
 wire \dpath.RF.R[10][0] ;
 wire \dpath.RF.R[10][10] ;
 wire \dpath.RF.R[10][11] ;
 wire \dpath.RF.R[10][12] ;
 wire \dpath.RF.R[10][13] ;
 wire \dpath.RF.R[10][14] ;
 wire \dpath.RF.R[10][15] ;
 wire \dpath.RF.R[10][16] ;
 wire \dpath.RF.R[10][17] ;
 wire \dpath.RF.R[10][18] ;
 wire \dpath.RF.R[10][19] ;
 wire \dpath.RF.R[10][1] ;
 wire \dpath.RF.R[10][20] ;
 wire \dpath.RF.R[10][21] ;
 wire \dpath.RF.R[10][22] ;
 wire \dpath.RF.R[10][23] ;
 wire \dpath.RF.R[10][24] ;
 wire \dpath.RF.R[10][25] ;
 wire \dpath.RF.R[10][26] ;
 wire \dpath.RF.R[10][27] ;
 wire \dpath.RF.R[10][28] ;
 wire \dpath.RF.R[10][29] ;
 wire \dpath.RF.R[10][2] ;
 wire \dpath.RF.R[10][30] ;
 wire \dpath.RF.R[10][31] ;
 wire \dpath.RF.R[10][3] ;
 wire \dpath.RF.R[10][4] ;
 wire \dpath.RF.R[10][5] ;
 wire \dpath.RF.R[10][6] ;
 wire \dpath.RF.R[10][7] ;
 wire \dpath.RF.R[10][8] ;
 wire \dpath.RF.R[10][9] ;
 wire \dpath.RF.R[11][0] ;
 wire \dpath.RF.R[11][10] ;
 wire \dpath.RF.R[11][11] ;
 wire \dpath.RF.R[11][12] ;
 wire \dpath.RF.R[11][13] ;
 wire \dpath.RF.R[11][14] ;
 wire \dpath.RF.R[11][15] ;
 wire \dpath.RF.R[11][16] ;
 wire \dpath.RF.R[11][17] ;
 wire \dpath.RF.R[11][18] ;
 wire \dpath.RF.R[11][19] ;
 wire \dpath.RF.R[11][1] ;
 wire \dpath.RF.R[11][20] ;
 wire \dpath.RF.R[11][21] ;
 wire \dpath.RF.R[11][22] ;
 wire \dpath.RF.R[11][23] ;
 wire \dpath.RF.R[11][24] ;
 wire \dpath.RF.R[11][25] ;
 wire \dpath.RF.R[11][26] ;
 wire \dpath.RF.R[11][27] ;
 wire \dpath.RF.R[11][28] ;
 wire \dpath.RF.R[11][29] ;
 wire \dpath.RF.R[11][2] ;
 wire \dpath.RF.R[11][30] ;
 wire \dpath.RF.R[11][31] ;
 wire \dpath.RF.R[11][3] ;
 wire \dpath.RF.R[11][4] ;
 wire \dpath.RF.R[11][5] ;
 wire \dpath.RF.R[11][6] ;
 wire \dpath.RF.R[11][7] ;
 wire \dpath.RF.R[11][8] ;
 wire \dpath.RF.R[11][9] ;
 wire \dpath.RF.R[12][0] ;
 wire \dpath.RF.R[12][10] ;
 wire \dpath.RF.R[12][11] ;
 wire \dpath.RF.R[12][12] ;
 wire \dpath.RF.R[12][13] ;
 wire \dpath.RF.R[12][14] ;
 wire \dpath.RF.R[12][15] ;
 wire \dpath.RF.R[12][16] ;
 wire \dpath.RF.R[12][17] ;
 wire \dpath.RF.R[12][18] ;
 wire \dpath.RF.R[12][19] ;
 wire \dpath.RF.R[12][1] ;
 wire \dpath.RF.R[12][20] ;
 wire \dpath.RF.R[12][21] ;
 wire \dpath.RF.R[12][22] ;
 wire \dpath.RF.R[12][23] ;
 wire \dpath.RF.R[12][24] ;
 wire \dpath.RF.R[12][25] ;
 wire \dpath.RF.R[12][26] ;
 wire \dpath.RF.R[12][27] ;
 wire \dpath.RF.R[12][28] ;
 wire \dpath.RF.R[12][29] ;
 wire \dpath.RF.R[12][2] ;
 wire \dpath.RF.R[12][30] ;
 wire \dpath.RF.R[12][31] ;
 wire \dpath.RF.R[12][3] ;
 wire \dpath.RF.R[12][4] ;
 wire \dpath.RF.R[12][5] ;
 wire \dpath.RF.R[12][6] ;
 wire \dpath.RF.R[12][7] ;
 wire \dpath.RF.R[12][8] ;
 wire \dpath.RF.R[12][9] ;
 wire \dpath.RF.R[13][0] ;
 wire \dpath.RF.R[13][10] ;
 wire \dpath.RF.R[13][11] ;
 wire \dpath.RF.R[13][12] ;
 wire \dpath.RF.R[13][13] ;
 wire \dpath.RF.R[13][14] ;
 wire \dpath.RF.R[13][15] ;
 wire \dpath.RF.R[13][16] ;
 wire \dpath.RF.R[13][17] ;
 wire \dpath.RF.R[13][18] ;
 wire \dpath.RF.R[13][19] ;
 wire \dpath.RF.R[13][1] ;
 wire \dpath.RF.R[13][20] ;
 wire \dpath.RF.R[13][21] ;
 wire \dpath.RF.R[13][22] ;
 wire \dpath.RF.R[13][23] ;
 wire \dpath.RF.R[13][24] ;
 wire \dpath.RF.R[13][25] ;
 wire \dpath.RF.R[13][26] ;
 wire \dpath.RF.R[13][27] ;
 wire \dpath.RF.R[13][28] ;
 wire \dpath.RF.R[13][29] ;
 wire \dpath.RF.R[13][2] ;
 wire \dpath.RF.R[13][30] ;
 wire \dpath.RF.R[13][31] ;
 wire \dpath.RF.R[13][3] ;
 wire \dpath.RF.R[13][4] ;
 wire \dpath.RF.R[13][5] ;
 wire \dpath.RF.R[13][6] ;
 wire \dpath.RF.R[13][7] ;
 wire \dpath.RF.R[13][8] ;
 wire \dpath.RF.R[13][9] ;
 wire \dpath.RF.R[14][0] ;
 wire \dpath.RF.R[14][10] ;
 wire \dpath.RF.R[14][11] ;
 wire \dpath.RF.R[14][12] ;
 wire \dpath.RF.R[14][13] ;
 wire \dpath.RF.R[14][14] ;
 wire \dpath.RF.R[14][15] ;
 wire \dpath.RF.R[14][16] ;
 wire \dpath.RF.R[14][17] ;
 wire \dpath.RF.R[14][18] ;
 wire \dpath.RF.R[14][19] ;
 wire \dpath.RF.R[14][1] ;
 wire \dpath.RF.R[14][20] ;
 wire \dpath.RF.R[14][21] ;
 wire \dpath.RF.R[14][22] ;
 wire \dpath.RF.R[14][23] ;
 wire \dpath.RF.R[14][24] ;
 wire \dpath.RF.R[14][25] ;
 wire \dpath.RF.R[14][26] ;
 wire \dpath.RF.R[14][27] ;
 wire \dpath.RF.R[14][28] ;
 wire \dpath.RF.R[14][29] ;
 wire \dpath.RF.R[14][2] ;
 wire \dpath.RF.R[14][30] ;
 wire \dpath.RF.R[14][31] ;
 wire \dpath.RF.R[14][3] ;
 wire \dpath.RF.R[14][4] ;
 wire \dpath.RF.R[14][5] ;
 wire \dpath.RF.R[14][6] ;
 wire \dpath.RF.R[14][7] ;
 wire \dpath.RF.R[14][8] ;
 wire \dpath.RF.R[14][9] ;
 wire \dpath.RF.R[15][0] ;
 wire \dpath.RF.R[15][10] ;
 wire \dpath.RF.R[15][11] ;
 wire \dpath.RF.R[15][12] ;
 wire \dpath.RF.R[15][13] ;
 wire \dpath.RF.R[15][14] ;
 wire \dpath.RF.R[15][15] ;
 wire \dpath.RF.R[15][16] ;
 wire \dpath.RF.R[15][17] ;
 wire \dpath.RF.R[15][18] ;
 wire \dpath.RF.R[15][19] ;
 wire \dpath.RF.R[15][1] ;
 wire \dpath.RF.R[15][20] ;
 wire \dpath.RF.R[15][21] ;
 wire \dpath.RF.R[15][22] ;
 wire \dpath.RF.R[15][23] ;
 wire \dpath.RF.R[15][24] ;
 wire \dpath.RF.R[15][25] ;
 wire \dpath.RF.R[15][26] ;
 wire \dpath.RF.R[15][27] ;
 wire \dpath.RF.R[15][28] ;
 wire \dpath.RF.R[15][29] ;
 wire \dpath.RF.R[15][2] ;
 wire \dpath.RF.R[15][30] ;
 wire \dpath.RF.R[15][31] ;
 wire \dpath.RF.R[15][3] ;
 wire \dpath.RF.R[15][4] ;
 wire \dpath.RF.R[15][5] ;
 wire \dpath.RF.R[15][6] ;
 wire \dpath.RF.R[15][7] ;
 wire \dpath.RF.R[15][8] ;
 wire \dpath.RF.R[15][9] ;
 wire \dpath.RF.R[16][0] ;
 wire \dpath.RF.R[16][10] ;
 wire \dpath.RF.R[16][11] ;
 wire \dpath.RF.R[16][12] ;
 wire \dpath.RF.R[16][13] ;
 wire \dpath.RF.R[16][14] ;
 wire \dpath.RF.R[16][15] ;
 wire \dpath.RF.R[16][16] ;
 wire \dpath.RF.R[16][17] ;
 wire \dpath.RF.R[16][18] ;
 wire \dpath.RF.R[16][19] ;
 wire \dpath.RF.R[16][1] ;
 wire \dpath.RF.R[16][20] ;
 wire \dpath.RF.R[16][21] ;
 wire \dpath.RF.R[16][22] ;
 wire \dpath.RF.R[16][23] ;
 wire \dpath.RF.R[16][24] ;
 wire \dpath.RF.R[16][25] ;
 wire \dpath.RF.R[16][26] ;
 wire \dpath.RF.R[16][27] ;
 wire \dpath.RF.R[16][28] ;
 wire \dpath.RF.R[16][29] ;
 wire \dpath.RF.R[16][2] ;
 wire \dpath.RF.R[16][30] ;
 wire \dpath.RF.R[16][31] ;
 wire \dpath.RF.R[16][3] ;
 wire \dpath.RF.R[16][4] ;
 wire \dpath.RF.R[16][5] ;
 wire \dpath.RF.R[16][6] ;
 wire \dpath.RF.R[16][7] ;
 wire \dpath.RF.R[16][8] ;
 wire \dpath.RF.R[16][9] ;
 wire \dpath.RF.R[17][0] ;
 wire \dpath.RF.R[17][10] ;
 wire \dpath.RF.R[17][11] ;
 wire \dpath.RF.R[17][12] ;
 wire \dpath.RF.R[17][13] ;
 wire \dpath.RF.R[17][14] ;
 wire \dpath.RF.R[17][15] ;
 wire \dpath.RF.R[17][16] ;
 wire \dpath.RF.R[17][17] ;
 wire \dpath.RF.R[17][18] ;
 wire \dpath.RF.R[17][19] ;
 wire \dpath.RF.R[17][1] ;
 wire \dpath.RF.R[17][20] ;
 wire \dpath.RF.R[17][21] ;
 wire \dpath.RF.R[17][22] ;
 wire \dpath.RF.R[17][23] ;
 wire \dpath.RF.R[17][24] ;
 wire \dpath.RF.R[17][25] ;
 wire \dpath.RF.R[17][26] ;
 wire \dpath.RF.R[17][27] ;
 wire \dpath.RF.R[17][28] ;
 wire \dpath.RF.R[17][29] ;
 wire \dpath.RF.R[17][2] ;
 wire \dpath.RF.R[17][30] ;
 wire \dpath.RF.R[17][31] ;
 wire \dpath.RF.R[17][3] ;
 wire \dpath.RF.R[17][4] ;
 wire \dpath.RF.R[17][5] ;
 wire \dpath.RF.R[17][6] ;
 wire \dpath.RF.R[17][7] ;
 wire \dpath.RF.R[17][8] ;
 wire \dpath.RF.R[17][9] ;
 wire \dpath.RF.R[18][0] ;
 wire \dpath.RF.R[18][10] ;
 wire \dpath.RF.R[18][11] ;
 wire \dpath.RF.R[18][12] ;
 wire \dpath.RF.R[18][13] ;
 wire \dpath.RF.R[18][14] ;
 wire \dpath.RF.R[18][15] ;
 wire \dpath.RF.R[18][16] ;
 wire \dpath.RF.R[18][17] ;
 wire \dpath.RF.R[18][18] ;
 wire \dpath.RF.R[18][19] ;
 wire \dpath.RF.R[18][1] ;
 wire \dpath.RF.R[18][20] ;
 wire \dpath.RF.R[18][21] ;
 wire \dpath.RF.R[18][22] ;
 wire \dpath.RF.R[18][23] ;
 wire \dpath.RF.R[18][24] ;
 wire \dpath.RF.R[18][25] ;
 wire \dpath.RF.R[18][26] ;
 wire \dpath.RF.R[18][27] ;
 wire \dpath.RF.R[18][28] ;
 wire \dpath.RF.R[18][29] ;
 wire \dpath.RF.R[18][2] ;
 wire \dpath.RF.R[18][30] ;
 wire \dpath.RF.R[18][31] ;
 wire \dpath.RF.R[18][3] ;
 wire \dpath.RF.R[18][4] ;
 wire \dpath.RF.R[18][5] ;
 wire \dpath.RF.R[18][6] ;
 wire \dpath.RF.R[18][7] ;
 wire \dpath.RF.R[18][8] ;
 wire \dpath.RF.R[18][9] ;
 wire \dpath.RF.R[19][0] ;
 wire \dpath.RF.R[19][10] ;
 wire \dpath.RF.R[19][11] ;
 wire \dpath.RF.R[19][12] ;
 wire \dpath.RF.R[19][13] ;
 wire \dpath.RF.R[19][14] ;
 wire \dpath.RF.R[19][15] ;
 wire \dpath.RF.R[19][16] ;
 wire \dpath.RF.R[19][17] ;
 wire \dpath.RF.R[19][18] ;
 wire \dpath.RF.R[19][19] ;
 wire \dpath.RF.R[19][1] ;
 wire \dpath.RF.R[19][20] ;
 wire \dpath.RF.R[19][21] ;
 wire \dpath.RF.R[19][22] ;
 wire \dpath.RF.R[19][23] ;
 wire \dpath.RF.R[19][24] ;
 wire \dpath.RF.R[19][25] ;
 wire \dpath.RF.R[19][26] ;
 wire \dpath.RF.R[19][27] ;
 wire \dpath.RF.R[19][28] ;
 wire \dpath.RF.R[19][29] ;
 wire \dpath.RF.R[19][2] ;
 wire \dpath.RF.R[19][30] ;
 wire \dpath.RF.R[19][31] ;
 wire \dpath.RF.R[19][3] ;
 wire \dpath.RF.R[19][4] ;
 wire \dpath.RF.R[19][5] ;
 wire \dpath.RF.R[19][6] ;
 wire \dpath.RF.R[19][7] ;
 wire \dpath.RF.R[19][8] ;
 wire \dpath.RF.R[19][9] ;
 wire \dpath.RF.R[1][0] ;
 wire \dpath.RF.R[1][10] ;
 wire \dpath.RF.R[1][11] ;
 wire \dpath.RF.R[1][12] ;
 wire \dpath.RF.R[1][13] ;
 wire \dpath.RF.R[1][14] ;
 wire \dpath.RF.R[1][15] ;
 wire \dpath.RF.R[1][16] ;
 wire \dpath.RF.R[1][17] ;
 wire \dpath.RF.R[1][18] ;
 wire \dpath.RF.R[1][19] ;
 wire \dpath.RF.R[1][1] ;
 wire \dpath.RF.R[1][20] ;
 wire \dpath.RF.R[1][21] ;
 wire \dpath.RF.R[1][22] ;
 wire \dpath.RF.R[1][23] ;
 wire \dpath.RF.R[1][24] ;
 wire \dpath.RF.R[1][25] ;
 wire \dpath.RF.R[1][26] ;
 wire \dpath.RF.R[1][27] ;
 wire \dpath.RF.R[1][28] ;
 wire \dpath.RF.R[1][29] ;
 wire \dpath.RF.R[1][2] ;
 wire \dpath.RF.R[1][30] ;
 wire \dpath.RF.R[1][31] ;
 wire \dpath.RF.R[1][3] ;
 wire \dpath.RF.R[1][4] ;
 wire \dpath.RF.R[1][5] ;
 wire \dpath.RF.R[1][6] ;
 wire \dpath.RF.R[1][7] ;
 wire \dpath.RF.R[1][8] ;
 wire \dpath.RF.R[1][9] ;
 wire \dpath.RF.R[20][0] ;
 wire \dpath.RF.R[20][10] ;
 wire \dpath.RF.R[20][11] ;
 wire \dpath.RF.R[20][12] ;
 wire \dpath.RF.R[20][13] ;
 wire \dpath.RF.R[20][14] ;
 wire \dpath.RF.R[20][15] ;
 wire \dpath.RF.R[20][16] ;
 wire \dpath.RF.R[20][17] ;
 wire \dpath.RF.R[20][18] ;
 wire \dpath.RF.R[20][19] ;
 wire \dpath.RF.R[20][1] ;
 wire \dpath.RF.R[20][20] ;
 wire \dpath.RF.R[20][21] ;
 wire \dpath.RF.R[20][22] ;
 wire \dpath.RF.R[20][23] ;
 wire \dpath.RF.R[20][24] ;
 wire \dpath.RF.R[20][25] ;
 wire \dpath.RF.R[20][26] ;
 wire \dpath.RF.R[20][27] ;
 wire \dpath.RF.R[20][28] ;
 wire \dpath.RF.R[20][29] ;
 wire \dpath.RF.R[20][2] ;
 wire \dpath.RF.R[20][30] ;
 wire \dpath.RF.R[20][31] ;
 wire \dpath.RF.R[20][3] ;
 wire \dpath.RF.R[20][4] ;
 wire \dpath.RF.R[20][5] ;
 wire \dpath.RF.R[20][6] ;
 wire \dpath.RF.R[20][7] ;
 wire \dpath.RF.R[20][8] ;
 wire \dpath.RF.R[20][9] ;
 wire \dpath.RF.R[21][0] ;
 wire \dpath.RF.R[21][10] ;
 wire \dpath.RF.R[21][11] ;
 wire \dpath.RF.R[21][12] ;
 wire \dpath.RF.R[21][13] ;
 wire \dpath.RF.R[21][14] ;
 wire \dpath.RF.R[21][15] ;
 wire \dpath.RF.R[21][16] ;
 wire \dpath.RF.R[21][17] ;
 wire \dpath.RF.R[21][18] ;
 wire \dpath.RF.R[21][19] ;
 wire \dpath.RF.R[21][1] ;
 wire \dpath.RF.R[21][20] ;
 wire \dpath.RF.R[21][21] ;
 wire \dpath.RF.R[21][22] ;
 wire \dpath.RF.R[21][23] ;
 wire \dpath.RF.R[21][24] ;
 wire \dpath.RF.R[21][25] ;
 wire \dpath.RF.R[21][26] ;
 wire \dpath.RF.R[21][27] ;
 wire \dpath.RF.R[21][28] ;
 wire \dpath.RF.R[21][29] ;
 wire \dpath.RF.R[21][2] ;
 wire \dpath.RF.R[21][30] ;
 wire \dpath.RF.R[21][31] ;
 wire \dpath.RF.R[21][3] ;
 wire \dpath.RF.R[21][4] ;
 wire \dpath.RF.R[21][5] ;
 wire \dpath.RF.R[21][6] ;
 wire \dpath.RF.R[21][7] ;
 wire \dpath.RF.R[21][8] ;
 wire \dpath.RF.R[21][9] ;
 wire \dpath.RF.R[22][0] ;
 wire \dpath.RF.R[22][10] ;
 wire \dpath.RF.R[22][11] ;
 wire \dpath.RF.R[22][12] ;
 wire \dpath.RF.R[22][13] ;
 wire \dpath.RF.R[22][14] ;
 wire \dpath.RF.R[22][15] ;
 wire \dpath.RF.R[22][16] ;
 wire \dpath.RF.R[22][17] ;
 wire \dpath.RF.R[22][18] ;
 wire \dpath.RF.R[22][19] ;
 wire \dpath.RF.R[22][1] ;
 wire \dpath.RF.R[22][20] ;
 wire \dpath.RF.R[22][21] ;
 wire \dpath.RF.R[22][22] ;
 wire \dpath.RF.R[22][23] ;
 wire \dpath.RF.R[22][24] ;
 wire \dpath.RF.R[22][25] ;
 wire \dpath.RF.R[22][26] ;
 wire \dpath.RF.R[22][27] ;
 wire \dpath.RF.R[22][28] ;
 wire \dpath.RF.R[22][29] ;
 wire \dpath.RF.R[22][2] ;
 wire \dpath.RF.R[22][30] ;
 wire \dpath.RF.R[22][31] ;
 wire \dpath.RF.R[22][3] ;
 wire \dpath.RF.R[22][4] ;
 wire \dpath.RF.R[22][5] ;
 wire \dpath.RF.R[22][6] ;
 wire \dpath.RF.R[22][7] ;
 wire \dpath.RF.R[22][8] ;
 wire \dpath.RF.R[22][9] ;
 wire \dpath.RF.R[23][0] ;
 wire \dpath.RF.R[23][10] ;
 wire \dpath.RF.R[23][11] ;
 wire \dpath.RF.R[23][12] ;
 wire \dpath.RF.R[23][13] ;
 wire \dpath.RF.R[23][14] ;
 wire \dpath.RF.R[23][15] ;
 wire \dpath.RF.R[23][16] ;
 wire \dpath.RF.R[23][17] ;
 wire \dpath.RF.R[23][18] ;
 wire \dpath.RF.R[23][19] ;
 wire \dpath.RF.R[23][1] ;
 wire \dpath.RF.R[23][20] ;
 wire \dpath.RF.R[23][21] ;
 wire \dpath.RF.R[23][22] ;
 wire \dpath.RF.R[23][23] ;
 wire \dpath.RF.R[23][24] ;
 wire \dpath.RF.R[23][25] ;
 wire \dpath.RF.R[23][26] ;
 wire \dpath.RF.R[23][27] ;
 wire \dpath.RF.R[23][28] ;
 wire \dpath.RF.R[23][29] ;
 wire \dpath.RF.R[23][2] ;
 wire \dpath.RF.R[23][30] ;
 wire \dpath.RF.R[23][31] ;
 wire \dpath.RF.R[23][3] ;
 wire \dpath.RF.R[23][4] ;
 wire \dpath.RF.R[23][5] ;
 wire \dpath.RF.R[23][6] ;
 wire \dpath.RF.R[23][7] ;
 wire \dpath.RF.R[23][8] ;
 wire \dpath.RF.R[23][9] ;
 wire \dpath.RF.R[24][0] ;
 wire \dpath.RF.R[24][10] ;
 wire \dpath.RF.R[24][11] ;
 wire \dpath.RF.R[24][12] ;
 wire \dpath.RF.R[24][13] ;
 wire \dpath.RF.R[24][14] ;
 wire \dpath.RF.R[24][15] ;
 wire \dpath.RF.R[24][16] ;
 wire \dpath.RF.R[24][17] ;
 wire \dpath.RF.R[24][18] ;
 wire \dpath.RF.R[24][19] ;
 wire \dpath.RF.R[24][1] ;
 wire \dpath.RF.R[24][20] ;
 wire \dpath.RF.R[24][21] ;
 wire \dpath.RF.R[24][22] ;
 wire \dpath.RF.R[24][23] ;
 wire \dpath.RF.R[24][24] ;
 wire \dpath.RF.R[24][25] ;
 wire \dpath.RF.R[24][26] ;
 wire \dpath.RF.R[24][27] ;
 wire \dpath.RF.R[24][28] ;
 wire \dpath.RF.R[24][29] ;
 wire \dpath.RF.R[24][2] ;
 wire \dpath.RF.R[24][30] ;
 wire \dpath.RF.R[24][31] ;
 wire \dpath.RF.R[24][3] ;
 wire \dpath.RF.R[24][4] ;
 wire \dpath.RF.R[24][5] ;
 wire \dpath.RF.R[24][6] ;
 wire \dpath.RF.R[24][7] ;
 wire \dpath.RF.R[24][8] ;
 wire \dpath.RF.R[24][9] ;
 wire \dpath.RF.R[25][0] ;
 wire \dpath.RF.R[25][10] ;
 wire \dpath.RF.R[25][11] ;
 wire \dpath.RF.R[25][12] ;
 wire \dpath.RF.R[25][13] ;
 wire \dpath.RF.R[25][14] ;
 wire \dpath.RF.R[25][15] ;
 wire \dpath.RF.R[25][16] ;
 wire \dpath.RF.R[25][17] ;
 wire \dpath.RF.R[25][18] ;
 wire \dpath.RF.R[25][19] ;
 wire \dpath.RF.R[25][1] ;
 wire \dpath.RF.R[25][20] ;
 wire \dpath.RF.R[25][21] ;
 wire \dpath.RF.R[25][22] ;
 wire \dpath.RF.R[25][23] ;
 wire \dpath.RF.R[25][24] ;
 wire \dpath.RF.R[25][25] ;
 wire \dpath.RF.R[25][26] ;
 wire \dpath.RF.R[25][27] ;
 wire \dpath.RF.R[25][28] ;
 wire \dpath.RF.R[25][29] ;
 wire \dpath.RF.R[25][2] ;
 wire \dpath.RF.R[25][30] ;
 wire \dpath.RF.R[25][31] ;
 wire \dpath.RF.R[25][3] ;
 wire \dpath.RF.R[25][4] ;
 wire \dpath.RF.R[25][5] ;
 wire \dpath.RF.R[25][6] ;
 wire \dpath.RF.R[25][7] ;
 wire \dpath.RF.R[25][8] ;
 wire \dpath.RF.R[25][9] ;
 wire \dpath.RF.R[26][0] ;
 wire \dpath.RF.R[26][10] ;
 wire \dpath.RF.R[26][11] ;
 wire \dpath.RF.R[26][12] ;
 wire \dpath.RF.R[26][13] ;
 wire \dpath.RF.R[26][14] ;
 wire \dpath.RF.R[26][15] ;
 wire \dpath.RF.R[26][16] ;
 wire \dpath.RF.R[26][17] ;
 wire \dpath.RF.R[26][18] ;
 wire \dpath.RF.R[26][19] ;
 wire \dpath.RF.R[26][1] ;
 wire \dpath.RF.R[26][20] ;
 wire \dpath.RF.R[26][21] ;
 wire \dpath.RF.R[26][22] ;
 wire \dpath.RF.R[26][23] ;
 wire \dpath.RF.R[26][24] ;
 wire \dpath.RF.R[26][25] ;
 wire \dpath.RF.R[26][26] ;
 wire \dpath.RF.R[26][27] ;
 wire \dpath.RF.R[26][28] ;
 wire \dpath.RF.R[26][29] ;
 wire \dpath.RF.R[26][2] ;
 wire \dpath.RF.R[26][30] ;
 wire \dpath.RF.R[26][31] ;
 wire \dpath.RF.R[26][3] ;
 wire \dpath.RF.R[26][4] ;
 wire \dpath.RF.R[26][5] ;
 wire \dpath.RF.R[26][6] ;
 wire \dpath.RF.R[26][7] ;
 wire \dpath.RF.R[26][8] ;
 wire \dpath.RF.R[26][9] ;
 wire \dpath.RF.R[27][0] ;
 wire \dpath.RF.R[27][10] ;
 wire \dpath.RF.R[27][11] ;
 wire \dpath.RF.R[27][12] ;
 wire \dpath.RF.R[27][13] ;
 wire \dpath.RF.R[27][14] ;
 wire \dpath.RF.R[27][15] ;
 wire \dpath.RF.R[27][16] ;
 wire \dpath.RF.R[27][17] ;
 wire \dpath.RF.R[27][18] ;
 wire \dpath.RF.R[27][19] ;
 wire \dpath.RF.R[27][1] ;
 wire \dpath.RF.R[27][20] ;
 wire \dpath.RF.R[27][21] ;
 wire \dpath.RF.R[27][22] ;
 wire \dpath.RF.R[27][23] ;
 wire \dpath.RF.R[27][24] ;
 wire \dpath.RF.R[27][25] ;
 wire \dpath.RF.R[27][26] ;
 wire \dpath.RF.R[27][27] ;
 wire \dpath.RF.R[27][28] ;
 wire \dpath.RF.R[27][29] ;
 wire \dpath.RF.R[27][2] ;
 wire \dpath.RF.R[27][30] ;
 wire \dpath.RF.R[27][31] ;
 wire \dpath.RF.R[27][3] ;
 wire \dpath.RF.R[27][4] ;
 wire \dpath.RF.R[27][5] ;
 wire \dpath.RF.R[27][6] ;
 wire \dpath.RF.R[27][7] ;
 wire \dpath.RF.R[27][8] ;
 wire \dpath.RF.R[27][9] ;
 wire \dpath.RF.R[28][0] ;
 wire \dpath.RF.R[28][10] ;
 wire \dpath.RF.R[28][11] ;
 wire \dpath.RF.R[28][12] ;
 wire \dpath.RF.R[28][13] ;
 wire \dpath.RF.R[28][14] ;
 wire \dpath.RF.R[28][15] ;
 wire \dpath.RF.R[28][16] ;
 wire \dpath.RF.R[28][17] ;
 wire \dpath.RF.R[28][18] ;
 wire \dpath.RF.R[28][19] ;
 wire \dpath.RF.R[28][1] ;
 wire \dpath.RF.R[28][20] ;
 wire \dpath.RF.R[28][21] ;
 wire \dpath.RF.R[28][22] ;
 wire \dpath.RF.R[28][23] ;
 wire \dpath.RF.R[28][24] ;
 wire \dpath.RF.R[28][25] ;
 wire \dpath.RF.R[28][26] ;
 wire \dpath.RF.R[28][27] ;
 wire \dpath.RF.R[28][28] ;
 wire \dpath.RF.R[28][29] ;
 wire \dpath.RF.R[28][2] ;
 wire \dpath.RF.R[28][30] ;
 wire \dpath.RF.R[28][31] ;
 wire \dpath.RF.R[28][3] ;
 wire \dpath.RF.R[28][4] ;
 wire \dpath.RF.R[28][5] ;
 wire \dpath.RF.R[28][6] ;
 wire \dpath.RF.R[28][7] ;
 wire \dpath.RF.R[28][8] ;
 wire \dpath.RF.R[28][9] ;
 wire \dpath.RF.R[29][0] ;
 wire \dpath.RF.R[29][10] ;
 wire \dpath.RF.R[29][11] ;
 wire \dpath.RF.R[29][12] ;
 wire \dpath.RF.R[29][13] ;
 wire \dpath.RF.R[29][14] ;
 wire \dpath.RF.R[29][15] ;
 wire \dpath.RF.R[29][16] ;
 wire \dpath.RF.R[29][17] ;
 wire \dpath.RF.R[29][18] ;
 wire \dpath.RF.R[29][19] ;
 wire \dpath.RF.R[29][1] ;
 wire \dpath.RF.R[29][20] ;
 wire \dpath.RF.R[29][21] ;
 wire \dpath.RF.R[29][22] ;
 wire \dpath.RF.R[29][23] ;
 wire \dpath.RF.R[29][24] ;
 wire \dpath.RF.R[29][25] ;
 wire \dpath.RF.R[29][26] ;
 wire \dpath.RF.R[29][27] ;
 wire \dpath.RF.R[29][28] ;
 wire \dpath.RF.R[29][29] ;
 wire \dpath.RF.R[29][2] ;
 wire \dpath.RF.R[29][30] ;
 wire \dpath.RF.R[29][31] ;
 wire \dpath.RF.R[29][3] ;
 wire \dpath.RF.R[29][4] ;
 wire \dpath.RF.R[29][5] ;
 wire \dpath.RF.R[29][6] ;
 wire \dpath.RF.R[29][7] ;
 wire \dpath.RF.R[29][8] ;
 wire \dpath.RF.R[29][9] ;
 wire \dpath.RF.R[2][0] ;
 wire \dpath.RF.R[2][10] ;
 wire \dpath.RF.R[2][11] ;
 wire \dpath.RF.R[2][12] ;
 wire \dpath.RF.R[2][13] ;
 wire \dpath.RF.R[2][14] ;
 wire \dpath.RF.R[2][15] ;
 wire \dpath.RF.R[2][16] ;
 wire \dpath.RF.R[2][17] ;
 wire \dpath.RF.R[2][18] ;
 wire \dpath.RF.R[2][19] ;
 wire \dpath.RF.R[2][1] ;
 wire \dpath.RF.R[2][20] ;
 wire \dpath.RF.R[2][21] ;
 wire \dpath.RF.R[2][22] ;
 wire \dpath.RF.R[2][23] ;
 wire \dpath.RF.R[2][24] ;
 wire \dpath.RF.R[2][25] ;
 wire \dpath.RF.R[2][26] ;
 wire \dpath.RF.R[2][27] ;
 wire \dpath.RF.R[2][28] ;
 wire \dpath.RF.R[2][29] ;
 wire \dpath.RF.R[2][2] ;
 wire \dpath.RF.R[2][30] ;
 wire \dpath.RF.R[2][31] ;
 wire \dpath.RF.R[2][3] ;
 wire \dpath.RF.R[2][4] ;
 wire \dpath.RF.R[2][5] ;
 wire \dpath.RF.R[2][6] ;
 wire \dpath.RF.R[2][7] ;
 wire \dpath.RF.R[2][8] ;
 wire \dpath.RF.R[2][9] ;
 wire \dpath.RF.R[30][0] ;
 wire \dpath.RF.R[30][10] ;
 wire \dpath.RF.R[30][11] ;
 wire \dpath.RF.R[30][12] ;
 wire \dpath.RF.R[30][13] ;
 wire \dpath.RF.R[30][14] ;
 wire \dpath.RF.R[30][15] ;
 wire \dpath.RF.R[30][16] ;
 wire \dpath.RF.R[30][17] ;
 wire \dpath.RF.R[30][18] ;
 wire \dpath.RF.R[30][19] ;
 wire \dpath.RF.R[30][1] ;
 wire \dpath.RF.R[30][20] ;
 wire \dpath.RF.R[30][21] ;
 wire \dpath.RF.R[30][22] ;
 wire \dpath.RF.R[30][23] ;
 wire \dpath.RF.R[30][24] ;
 wire \dpath.RF.R[30][25] ;
 wire \dpath.RF.R[30][26] ;
 wire \dpath.RF.R[30][27] ;
 wire \dpath.RF.R[30][28] ;
 wire \dpath.RF.R[30][29] ;
 wire \dpath.RF.R[30][2] ;
 wire \dpath.RF.R[30][30] ;
 wire \dpath.RF.R[30][31] ;
 wire \dpath.RF.R[30][3] ;
 wire \dpath.RF.R[30][4] ;
 wire \dpath.RF.R[30][5] ;
 wire \dpath.RF.R[30][6] ;
 wire \dpath.RF.R[30][7] ;
 wire \dpath.RF.R[30][8] ;
 wire \dpath.RF.R[30][9] ;
 wire \dpath.RF.R[31][0] ;
 wire \dpath.RF.R[31][10] ;
 wire \dpath.RF.R[31][11] ;
 wire \dpath.RF.R[31][12] ;
 wire \dpath.RF.R[31][13] ;
 wire \dpath.RF.R[31][14] ;
 wire \dpath.RF.R[31][15] ;
 wire \dpath.RF.R[31][16] ;
 wire \dpath.RF.R[31][17] ;
 wire \dpath.RF.R[31][18] ;
 wire \dpath.RF.R[31][19] ;
 wire \dpath.RF.R[31][1] ;
 wire \dpath.RF.R[31][20] ;
 wire \dpath.RF.R[31][21] ;
 wire \dpath.RF.R[31][22] ;
 wire \dpath.RF.R[31][23] ;
 wire \dpath.RF.R[31][24] ;
 wire \dpath.RF.R[31][25] ;
 wire \dpath.RF.R[31][26] ;
 wire \dpath.RF.R[31][27] ;
 wire \dpath.RF.R[31][28] ;
 wire \dpath.RF.R[31][29] ;
 wire \dpath.RF.R[31][2] ;
 wire \dpath.RF.R[31][30] ;
 wire \dpath.RF.R[31][31] ;
 wire \dpath.RF.R[31][3] ;
 wire \dpath.RF.R[31][4] ;
 wire \dpath.RF.R[31][5] ;
 wire \dpath.RF.R[31][6] ;
 wire \dpath.RF.R[31][7] ;
 wire \dpath.RF.R[31][8] ;
 wire \dpath.RF.R[31][9] ;
 wire \dpath.RF.R[3][0] ;
 wire \dpath.RF.R[3][10] ;
 wire \dpath.RF.R[3][11] ;
 wire \dpath.RF.R[3][12] ;
 wire \dpath.RF.R[3][13] ;
 wire \dpath.RF.R[3][14] ;
 wire \dpath.RF.R[3][15] ;
 wire \dpath.RF.R[3][16] ;
 wire \dpath.RF.R[3][17] ;
 wire \dpath.RF.R[3][18] ;
 wire \dpath.RF.R[3][19] ;
 wire \dpath.RF.R[3][1] ;
 wire \dpath.RF.R[3][20] ;
 wire \dpath.RF.R[3][21] ;
 wire \dpath.RF.R[3][22] ;
 wire \dpath.RF.R[3][23] ;
 wire \dpath.RF.R[3][24] ;
 wire \dpath.RF.R[3][25] ;
 wire \dpath.RF.R[3][26] ;
 wire \dpath.RF.R[3][27] ;
 wire \dpath.RF.R[3][28] ;
 wire \dpath.RF.R[3][29] ;
 wire \dpath.RF.R[3][2] ;
 wire \dpath.RF.R[3][30] ;
 wire \dpath.RF.R[3][31] ;
 wire \dpath.RF.R[3][3] ;
 wire \dpath.RF.R[3][4] ;
 wire \dpath.RF.R[3][5] ;
 wire \dpath.RF.R[3][6] ;
 wire \dpath.RF.R[3][7] ;
 wire \dpath.RF.R[3][8] ;
 wire \dpath.RF.R[3][9] ;
 wire \dpath.RF.R[4][0] ;
 wire \dpath.RF.R[4][10] ;
 wire \dpath.RF.R[4][11] ;
 wire \dpath.RF.R[4][12] ;
 wire \dpath.RF.R[4][13] ;
 wire \dpath.RF.R[4][14] ;
 wire \dpath.RF.R[4][15] ;
 wire \dpath.RF.R[4][16] ;
 wire \dpath.RF.R[4][17] ;
 wire \dpath.RF.R[4][18] ;
 wire \dpath.RF.R[4][19] ;
 wire \dpath.RF.R[4][1] ;
 wire \dpath.RF.R[4][20] ;
 wire \dpath.RF.R[4][21] ;
 wire \dpath.RF.R[4][22] ;
 wire \dpath.RF.R[4][23] ;
 wire \dpath.RF.R[4][24] ;
 wire \dpath.RF.R[4][25] ;
 wire \dpath.RF.R[4][26] ;
 wire \dpath.RF.R[4][27] ;
 wire \dpath.RF.R[4][28] ;
 wire \dpath.RF.R[4][29] ;
 wire \dpath.RF.R[4][2] ;
 wire \dpath.RF.R[4][30] ;
 wire \dpath.RF.R[4][31] ;
 wire \dpath.RF.R[4][3] ;
 wire \dpath.RF.R[4][4] ;
 wire \dpath.RF.R[4][5] ;
 wire \dpath.RF.R[4][6] ;
 wire \dpath.RF.R[4][7] ;
 wire \dpath.RF.R[4][8] ;
 wire \dpath.RF.R[4][9] ;
 wire \dpath.RF.R[5][0] ;
 wire \dpath.RF.R[5][10] ;
 wire \dpath.RF.R[5][11] ;
 wire \dpath.RF.R[5][12] ;
 wire \dpath.RF.R[5][13] ;
 wire \dpath.RF.R[5][14] ;
 wire \dpath.RF.R[5][15] ;
 wire \dpath.RF.R[5][16] ;
 wire \dpath.RF.R[5][17] ;
 wire \dpath.RF.R[5][18] ;
 wire \dpath.RF.R[5][19] ;
 wire \dpath.RF.R[5][1] ;
 wire \dpath.RF.R[5][20] ;
 wire \dpath.RF.R[5][21] ;
 wire \dpath.RF.R[5][22] ;
 wire \dpath.RF.R[5][23] ;
 wire \dpath.RF.R[5][24] ;
 wire \dpath.RF.R[5][25] ;
 wire \dpath.RF.R[5][26] ;
 wire \dpath.RF.R[5][27] ;
 wire \dpath.RF.R[5][28] ;
 wire \dpath.RF.R[5][29] ;
 wire \dpath.RF.R[5][2] ;
 wire \dpath.RF.R[5][30] ;
 wire \dpath.RF.R[5][31] ;
 wire \dpath.RF.R[5][3] ;
 wire \dpath.RF.R[5][4] ;
 wire \dpath.RF.R[5][5] ;
 wire \dpath.RF.R[5][6] ;
 wire \dpath.RF.R[5][7] ;
 wire \dpath.RF.R[5][8] ;
 wire \dpath.RF.R[5][9] ;
 wire \dpath.RF.R[6][0] ;
 wire \dpath.RF.R[6][10] ;
 wire \dpath.RF.R[6][11] ;
 wire \dpath.RF.R[6][12] ;
 wire \dpath.RF.R[6][13] ;
 wire \dpath.RF.R[6][14] ;
 wire \dpath.RF.R[6][15] ;
 wire \dpath.RF.R[6][16] ;
 wire \dpath.RF.R[6][17] ;
 wire \dpath.RF.R[6][18] ;
 wire \dpath.RF.R[6][19] ;
 wire \dpath.RF.R[6][1] ;
 wire \dpath.RF.R[6][20] ;
 wire \dpath.RF.R[6][21] ;
 wire \dpath.RF.R[6][22] ;
 wire \dpath.RF.R[6][23] ;
 wire \dpath.RF.R[6][24] ;
 wire \dpath.RF.R[6][25] ;
 wire \dpath.RF.R[6][26] ;
 wire \dpath.RF.R[6][27] ;
 wire \dpath.RF.R[6][28] ;
 wire \dpath.RF.R[6][29] ;
 wire \dpath.RF.R[6][2] ;
 wire \dpath.RF.R[6][30] ;
 wire \dpath.RF.R[6][31] ;
 wire \dpath.RF.R[6][3] ;
 wire \dpath.RF.R[6][4] ;
 wire \dpath.RF.R[6][5] ;
 wire \dpath.RF.R[6][6] ;
 wire \dpath.RF.R[6][7] ;
 wire \dpath.RF.R[6][8] ;
 wire \dpath.RF.R[6][9] ;
 wire \dpath.RF.R[7][0] ;
 wire \dpath.RF.R[7][10] ;
 wire \dpath.RF.R[7][11] ;
 wire \dpath.RF.R[7][12] ;
 wire \dpath.RF.R[7][13] ;
 wire \dpath.RF.R[7][14] ;
 wire \dpath.RF.R[7][15] ;
 wire \dpath.RF.R[7][16] ;
 wire \dpath.RF.R[7][17] ;
 wire \dpath.RF.R[7][18] ;
 wire \dpath.RF.R[7][19] ;
 wire \dpath.RF.R[7][1] ;
 wire \dpath.RF.R[7][20] ;
 wire \dpath.RF.R[7][21] ;
 wire \dpath.RF.R[7][22] ;
 wire \dpath.RF.R[7][23] ;
 wire \dpath.RF.R[7][24] ;
 wire \dpath.RF.R[7][25] ;
 wire \dpath.RF.R[7][26] ;
 wire \dpath.RF.R[7][27] ;
 wire \dpath.RF.R[7][28] ;
 wire \dpath.RF.R[7][29] ;
 wire \dpath.RF.R[7][2] ;
 wire \dpath.RF.R[7][30] ;
 wire \dpath.RF.R[7][31] ;
 wire \dpath.RF.R[7][3] ;
 wire \dpath.RF.R[7][4] ;
 wire \dpath.RF.R[7][5] ;
 wire \dpath.RF.R[7][6] ;
 wire \dpath.RF.R[7][7] ;
 wire \dpath.RF.R[7][8] ;
 wire \dpath.RF.R[7][9] ;
 wire \dpath.RF.R[8][0] ;
 wire \dpath.RF.R[8][10] ;
 wire \dpath.RF.R[8][11] ;
 wire \dpath.RF.R[8][12] ;
 wire \dpath.RF.R[8][13] ;
 wire \dpath.RF.R[8][14] ;
 wire \dpath.RF.R[8][15] ;
 wire \dpath.RF.R[8][16] ;
 wire \dpath.RF.R[8][17] ;
 wire \dpath.RF.R[8][18] ;
 wire \dpath.RF.R[8][19] ;
 wire \dpath.RF.R[8][1] ;
 wire \dpath.RF.R[8][20] ;
 wire \dpath.RF.R[8][21] ;
 wire \dpath.RF.R[8][22] ;
 wire \dpath.RF.R[8][23] ;
 wire \dpath.RF.R[8][24] ;
 wire \dpath.RF.R[8][25] ;
 wire \dpath.RF.R[8][26] ;
 wire \dpath.RF.R[8][27] ;
 wire \dpath.RF.R[8][28] ;
 wire \dpath.RF.R[8][29] ;
 wire \dpath.RF.R[8][2] ;
 wire \dpath.RF.R[8][30] ;
 wire \dpath.RF.R[8][31] ;
 wire \dpath.RF.R[8][3] ;
 wire \dpath.RF.R[8][4] ;
 wire \dpath.RF.R[8][5] ;
 wire \dpath.RF.R[8][6] ;
 wire \dpath.RF.R[8][7] ;
 wire \dpath.RF.R[8][8] ;
 wire \dpath.RF.R[8][9] ;
 wire \dpath.RF.R[9][0] ;
 wire \dpath.RF.R[9][10] ;
 wire \dpath.RF.R[9][11] ;
 wire \dpath.RF.R[9][12] ;
 wire \dpath.RF.R[9][13] ;
 wire \dpath.RF.R[9][14] ;
 wire \dpath.RF.R[9][15] ;
 wire \dpath.RF.R[9][16] ;
 wire \dpath.RF.R[9][17] ;
 wire \dpath.RF.R[9][18] ;
 wire \dpath.RF.R[9][19] ;
 wire \dpath.RF.R[9][1] ;
 wire \dpath.RF.R[9][20] ;
 wire \dpath.RF.R[9][21] ;
 wire \dpath.RF.R[9][22] ;
 wire \dpath.RF.R[9][23] ;
 wire \dpath.RF.R[9][24] ;
 wire \dpath.RF.R[9][25] ;
 wire \dpath.RF.R[9][26] ;
 wire \dpath.RF.R[9][27] ;
 wire \dpath.RF.R[9][28] ;
 wire \dpath.RF.R[9][29] ;
 wire \dpath.RF.R[9][2] ;
 wire \dpath.RF.R[9][30] ;
 wire \dpath.RF.R[9][31] ;
 wire \dpath.RF.R[9][3] ;
 wire \dpath.RF.R[9][4] ;
 wire \dpath.RF.R[9][5] ;
 wire \dpath.RF.R[9][6] ;
 wire \dpath.RF.R[9][7] ;
 wire \dpath.RF.R[9][8] ;
 wire \dpath.RF.R[9][9] ;
 wire \dpath.RF.wdata[0] ;
 wire \dpath.RF.wdata[10] ;
 wire \dpath.RF.wdata[11] ;
 wire \dpath.RF.wdata[12] ;
 wire \dpath.RF.wdata[13] ;
 wire \dpath.RF.wdata[14] ;
 wire \dpath.RF.wdata[15] ;
 wire \dpath.RF.wdata[16] ;
 wire \dpath.RF.wdata[17] ;
 wire \dpath.RF.wdata[18] ;
 wire \dpath.RF.wdata[19] ;
 wire \dpath.RF.wdata[1] ;
 wire \dpath.RF.wdata[20] ;
 wire \dpath.RF.wdata[21] ;
 wire \dpath.RF.wdata[22] ;
 wire \dpath.RF.wdata[23] ;
 wire \dpath.RF.wdata[24] ;
 wire \dpath.RF.wdata[25] ;
 wire \dpath.RF.wdata[26] ;
 wire \dpath.RF.wdata[27] ;
 wire \dpath.RF.wdata[28] ;
 wire \dpath.RF.wdata[29] ;
 wire \dpath.RF.wdata[2] ;
 wire \dpath.RF.wdata[30] ;
 wire \dpath.RF.wdata[31] ;
 wire \dpath.RF.wdata[3] ;
 wire \dpath.RF.wdata[4] ;
 wire \dpath.RF.wdata[5] ;
 wire \dpath.RF.wdata[6] ;
 wire \dpath.RF.wdata[7] ;
 wire \dpath.RF.wdata[8] ;
 wire \dpath.RF.wdata[9] ;
 wire \dpath.alu.adder.in0[0] ;
 wire \dpath.alu.adder.in0[10] ;
 wire \dpath.alu.adder.in0[11] ;
 wire \dpath.alu.adder.in0[12] ;
 wire \dpath.alu.adder.in0[13] ;
 wire \dpath.alu.adder.in0[14] ;
 wire \dpath.alu.adder.in0[15] ;
 wire \dpath.alu.adder.in0[16] ;
 wire \dpath.alu.adder.in0[17] ;
 wire \dpath.alu.adder.in0[18] ;
 wire \dpath.alu.adder.in0[19] ;
 wire \dpath.alu.adder.in0[1] ;
 wire \dpath.alu.adder.in0[20] ;
 wire \dpath.alu.adder.in0[21] ;
 wire \dpath.alu.adder.in0[22] ;
 wire \dpath.alu.adder.in0[23] ;
 wire \dpath.alu.adder.in0[24] ;
 wire \dpath.alu.adder.in0[25] ;
 wire \dpath.alu.adder.in0[26] ;
 wire \dpath.alu.adder.in0[27] ;
 wire \dpath.alu.adder.in0[28] ;
 wire \dpath.alu.adder.in0[29] ;
 wire \dpath.alu.adder.in0[2] ;
 wire \dpath.alu.adder.in0[30] ;
 wire \dpath.alu.adder.in0[31] ;
 wire \dpath.alu.adder.in0[3] ;
 wire \dpath.alu.adder.in0[4] ;
 wire \dpath.alu.adder.in0[5] ;
 wire \dpath.alu.adder.in0[6] ;
 wire \dpath.alu.adder.in0[7] ;
 wire \dpath.alu.adder.in0[8] ;
 wire \dpath.alu.adder.in0[9] ;
 wire \dpath.alu.adder.in1[0] ;
 wire \dpath.alu.adder.in1[10] ;
 wire \dpath.alu.adder.in1[11] ;
 wire \dpath.alu.adder.in1[12] ;
 wire \dpath.alu.adder.in1[13] ;
 wire \dpath.alu.adder.in1[14] ;
 wire \dpath.alu.adder.in1[15] ;
 wire \dpath.alu.adder.in1[16] ;
 wire \dpath.alu.adder.in1[17] ;
 wire \dpath.alu.adder.in1[18] ;
 wire \dpath.alu.adder.in1[19] ;
 wire \dpath.alu.adder.in1[1] ;
 wire \dpath.alu.adder.in1[20] ;
 wire \dpath.alu.adder.in1[21] ;
 wire \dpath.alu.adder.in1[22] ;
 wire \dpath.alu.adder.in1[23] ;
 wire \dpath.alu.adder.in1[24] ;
 wire \dpath.alu.adder.in1[25] ;
 wire \dpath.alu.adder.in1[26] ;
 wire \dpath.alu.adder.in1[27] ;
 wire \dpath.alu.adder.in1[28] ;
 wire \dpath.alu.adder.in1[29] ;
 wire \dpath.alu.adder.in1[2] ;
 wire \dpath.alu.adder.in1[30] ;
 wire \dpath.alu.adder.in1[31] ;
 wire \dpath.alu.adder.in1[3] ;
 wire \dpath.alu.adder.in1[4] ;
 wire \dpath.alu.adder.in1[5] ;
 wire \dpath.alu.adder.in1[6] ;
 wire \dpath.alu.adder.in1[7] ;
 wire \dpath.alu.adder.in1[8] ;
 wire \dpath.alu.adder.in1[9] ;
 wire \dpath.btarg_DX.q[0] ;
 wire \dpath.btarg_DX.q[10] ;
 wire \dpath.btarg_DX.q[11] ;
 wire \dpath.btarg_DX.q[12] ;
 wire \dpath.btarg_DX.q[13] ;
 wire \dpath.btarg_DX.q[14] ;
 wire \dpath.btarg_DX.q[15] ;
 wire \dpath.btarg_DX.q[16] ;
 wire \dpath.btarg_DX.q[17] ;
 wire \dpath.btarg_DX.q[18] ;
 wire \dpath.btarg_DX.q[19] ;
 wire \dpath.btarg_DX.q[1] ;
 wire \dpath.btarg_DX.q[20] ;
 wire \dpath.btarg_DX.q[21] ;
 wire \dpath.btarg_DX.q[22] ;
 wire \dpath.btarg_DX.q[23] ;
 wire \dpath.btarg_DX.q[24] ;
 wire \dpath.btarg_DX.q[25] ;
 wire \dpath.btarg_DX.q[26] ;
 wire \dpath.btarg_DX.q[27] ;
 wire \dpath.btarg_DX.q[28] ;
 wire \dpath.btarg_DX.q[29] ;
 wire \dpath.btarg_DX.q[2] ;
 wire \dpath.btarg_DX.q[30] ;
 wire \dpath.btarg_DX.q[31] ;
 wire \dpath.btarg_DX.q[3] ;
 wire \dpath.btarg_DX.q[4] ;
 wire \dpath.btarg_DX.q[5] ;
 wire \dpath.btarg_DX.q[6] ;
 wire \dpath.btarg_DX.q[7] ;
 wire \dpath.btarg_DX.q[8] ;
 wire \dpath.btarg_DX.q[9] ;
 wire \dpath.csrr[0] ;
 wire \dpath.csrr[10] ;
 wire \dpath.csrr[11] ;
 wire \dpath.csrr[12] ;
 wire \dpath.csrr[13] ;
 wire \dpath.csrr[14] ;
 wire \dpath.csrr[15] ;
 wire \dpath.csrr[16] ;
 wire \dpath.csrr[17] ;
 wire \dpath.csrr[18] ;
 wire \dpath.csrr[19] ;
 wire \dpath.csrr[1] ;
 wire \dpath.csrr[20] ;
 wire \dpath.csrr[21] ;
 wire \dpath.csrr[22] ;
 wire \dpath.csrr[23] ;
 wire \dpath.csrr[24] ;
 wire \dpath.csrr[25] ;
 wire \dpath.csrr[26] ;
 wire \dpath.csrr[27] ;
 wire \dpath.csrr[28] ;
 wire \dpath.csrr[29] ;
 wire \dpath.csrr[2] ;
 wire \dpath.csrr[30] ;
 wire \dpath.csrr[31] ;
 wire \dpath.csrr[3] ;
 wire \dpath.csrr[4] ;
 wire \dpath.csrr[5] ;
 wire \dpath.csrr[6] ;
 wire \dpath.csrr[7] ;
 wire \dpath.csrr[8] ;
 wire \dpath.csrr[9] ;
 wire \dpath.csrw_out0.d[0] ;
 wire \dpath.csrw_out0.d[10] ;
 wire \dpath.csrw_out0.d[11] ;
 wire \dpath.csrw_out0.d[12] ;
 wire \dpath.csrw_out0.d[13] ;
 wire \dpath.csrw_out0.d[14] ;
 wire \dpath.csrw_out0.d[15] ;
 wire \dpath.csrw_out0.d[16] ;
 wire \dpath.csrw_out0.d[17] ;
 wire \dpath.csrw_out0.d[18] ;
 wire \dpath.csrw_out0.d[19] ;
 wire \dpath.csrw_out0.d[1] ;
 wire \dpath.csrw_out0.d[20] ;
 wire \dpath.csrw_out0.d[21] ;
 wire \dpath.csrw_out0.d[22] ;
 wire \dpath.csrw_out0.d[23] ;
 wire \dpath.csrw_out0.d[24] ;
 wire \dpath.csrw_out0.d[25] ;
 wire \dpath.csrw_out0.d[26] ;
 wire \dpath.csrw_out0.d[27] ;
 wire \dpath.csrw_out0.d[28] ;
 wire \dpath.csrw_out0.d[29] ;
 wire \dpath.csrw_out0.d[2] ;
 wire \dpath.csrw_out0.d[30] ;
 wire \dpath.csrw_out0.d[31] ;
 wire \dpath.csrw_out0.d[3] ;
 wire \dpath.csrw_out0.d[4] ;
 wire \dpath.csrw_out0.d[5] ;
 wire \dpath.csrw_out0.d[6] ;
 wire \dpath.csrw_out0.d[7] ;
 wire \dpath.csrw_out0.d[8] ;
 wire \dpath.csrw_out0.d[9] ;
 wire \dpath.csrw_out_DX.q[0] ;
 wire \dpath.csrw_out_DX.q[10] ;
 wire \dpath.csrw_out_DX.q[11] ;
 wire \dpath.csrw_out_DX.q[12] ;
 wire \dpath.csrw_out_DX.q[13] ;
 wire \dpath.csrw_out_DX.q[14] ;
 wire \dpath.csrw_out_DX.q[15] ;
 wire \dpath.csrw_out_DX.q[16] ;
 wire \dpath.csrw_out_DX.q[17] ;
 wire \dpath.csrw_out_DX.q[18] ;
 wire \dpath.csrw_out_DX.q[19] ;
 wire \dpath.csrw_out_DX.q[1] ;
 wire \dpath.csrw_out_DX.q[20] ;
 wire \dpath.csrw_out_DX.q[21] ;
 wire \dpath.csrw_out_DX.q[22] ;
 wire \dpath.csrw_out_DX.q[23] ;
 wire \dpath.csrw_out_DX.q[24] ;
 wire \dpath.csrw_out_DX.q[25] ;
 wire \dpath.csrw_out_DX.q[26] ;
 wire \dpath.csrw_out_DX.q[27] ;
 wire \dpath.csrw_out_DX.q[28] ;
 wire \dpath.csrw_out_DX.q[29] ;
 wire \dpath.csrw_out_DX.q[2] ;
 wire \dpath.csrw_out_DX.q[30] ;
 wire \dpath.csrw_out_DX.q[31] ;
 wire \dpath.csrw_out_DX.q[3] ;
 wire \dpath.csrw_out_DX.q[4] ;
 wire \dpath.csrw_out_DX.q[5] ;
 wire \dpath.csrw_out_DX.q[6] ;
 wire \dpath.csrw_out_DX.q[7] ;
 wire \dpath.csrw_out_DX.q[8] ;
 wire \dpath.csrw_out_DX.q[9] ;
 wire \dpath.csrw_out_MW.d[0] ;
 wire \dpath.csrw_out_MW.d[10] ;
 wire \dpath.csrw_out_MW.d[11] ;
 wire \dpath.csrw_out_MW.d[12] ;
 wire \dpath.csrw_out_MW.d[13] ;
 wire \dpath.csrw_out_MW.d[14] ;
 wire \dpath.csrw_out_MW.d[15] ;
 wire \dpath.csrw_out_MW.d[16] ;
 wire \dpath.csrw_out_MW.d[17] ;
 wire \dpath.csrw_out_MW.d[18] ;
 wire \dpath.csrw_out_MW.d[19] ;
 wire \dpath.csrw_out_MW.d[1] ;
 wire \dpath.csrw_out_MW.d[20] ;
 wire \dpath.csrw_out_MW.d[21] ;
 wire \dpath.csrw_out_MW.d[22] ;
 wire \dpath.csrw_out_MW.d[23] ;
 wire \dpath.csrw_out_MW.d[24] ;
 wire \dpath.csrw_out_MW.d[25] ;
 wire \dpath.csrw_out_MW.d[26] ;
 wire \dpath.csrw_out_MW.d[27] ;
 wire \dpath.csrw_out_MW.d[28] ;
 wire \dpath.csrw_out_MW.d[29] ;
 wire \dpath.csrw_out_MW.d[2] ;
 wire \dpath.csrw_out_MW.d[30] ;
 wire \dpath.csrw_out_MW.d[31] ;
 wire \dpath.csrw_out_MW.d[3] ;
 wire \dpath.csrw_out_MW.d[4] ;
 wire \dpath.csrw_out_MW.d[5] ;
 wire \dpath.csrw_out_MW.d[6] ;
 wire \dpath.csrw_out_MW.d[7] ;
 wire \dpath.csrw_out_MW.d[8] ;
 wire \dpath.csrw_out_MW.d[9] ;
 wire \dpath.inst_pc[0] ;
 wire \dpath.inst_pc[10] ;
 wire \dpath.inst_pc[11] ;
 wire \dpath.inst_pc[12] ;
 wire \dpath.inst_pc[13] ;
 wire \dpath.inst_pc[14] ;
 wire \dpath.inst_pc[15] ;
 wire \dpath.inst_pc[16] ;
 wire \dpath.inst_pc[17] ;
 wire \dpath.inst_pc[18] ;
 wire \dpath.inst_pc[19] ;
 wire \dpath.inst_pc[1] ;
 wire \dpath.inst_pc[20] ;
 wire \dpath.inst_pc[21] ;
 wire \dpath.inst_pc[22] ;
 wire \dpath.inst_pc[23] ;
 wire \dpath.inst_pc[24] ;
 wire \dpath.inst_pc[25] ;
 wire \dpath.inst_pc[26] ;
 wire \dpath.inst_pc[27] ;
 wire \dpath.inst_pc[28] ;
 wire \dpath.inst_pc[29] ;
 wire \dpath.inst_pc[2] ;
 wire \dpath.inst_pc[30] ;
 wire \dpath.inst_pc[31] ;
 wire \dpath.inst_pc[3] ;
 wire \dpath.inst_pc[4] ;
 wire \dpath.inst_pc[5] ;
 wire \dpath.inst_pc[6] ;
 wire \dpath.inst_pc[7] ;
 wire \dpath.inst_pc[8] ;
 wire \dpath.inst_pc[9] ;
 wire \dpath.sd_DX.q[0] ;
 wire \dpath.sd_DX.q[10] ;
 wire \dpath.sd_DX.q[11] ;
 wire \dpath.sd_DX.q[12] ;
 wire \dpath.sd_DX.q[13] ;
 wire \dpath.sd_DX.q[14] ;
 wire \dpath.sd_DX.q[15] ;
 wire \dpath.sd_DX.q[16] ;
 wire \dpath.sd_DX.q[17] ;
 wire \dpath.sd_DX.q[18] ;
 wire \dpath.sd_DX.q[19] ;
 wire \dpath.sd_DX.q[1] ;
 wire \dpath.sd_DX.q[20] ;
 wire \dpath.sd_DX.q[21] ;
 wire \dpath.sd_DX.q[22] ;
 wire \dpath.sd_DX.q[23] ;
 wire \dpath.sd_DX.q[24] ;
 wire \dpath.sd_DX.q[25] ;
 wire \dpath.sd_DX.q[26] ;
 wire \dpath.sd_DX.q[27] ;
 wire \dpath.sd_DX.q[28] ;
 wire \dpath.sd_DX.q[29] ;
 wire \dpath.sd_DX.q[2] ;
 wire \dpath.sd_DX.q[30] ;
 wire \dpath.sd_DX.q[31] ;
 wire \dpath.sd_DX.q[3] ;
 wire \dpath.sd_DX.q[4] ;
 wire \dpath.sd_DX.q[5] ;
 wire \dpath.sd_DX.q[6] ;
 wire \dpath.sd_DX.q[7] ;
 wire \dpath.sd_DX.q[8] ;
 wire \dpath.sd_DX.q[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net303;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net317;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net342;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net356;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net358;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net363;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net368;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net371;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net372;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net373;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net374;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net375;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net376;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_01421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_01421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_01421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_01421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\dpath.sd_DX.q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_01219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(_06022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(_06022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_01140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_01140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_01140_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_01225_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_01225_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_01225_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_01417_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_01944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_05989_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\dpath.sd_DX.q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net3359));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__A (.DIODE(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__A (.DIODE(\ctrl.d2c_inst[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__A (.DIODE(\ctrl.d2c_inst[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B1 (.DIODE(_01804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__S (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__S (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__S (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__S (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__S (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__S (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__A0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A0 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__S (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A0 (.DIODE(\dpath.RF.wdata[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__S (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__A0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__A0 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__S (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__S (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__A0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__S (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__S (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__S (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__S (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__A (.DIODE(\dpath.alu.adder.in0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__A (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A (.DIODE(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__B (.DIODE(\dpath.alu.adder.in1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A (.DIODE(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B (.DIODE(\dpath.alu.adder.in1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__B (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__B (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A (.DIODE(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__B (.DIODE(\dpath.alu.adder.in1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A (.DIODE(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B (.DIODE(\dpath.alu.adder.in1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__B (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__B (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__B (.DIODE(\dpath.alu.adder.in1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B (.DIODE(\dpath.alu.adder.in1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(\dpath.alu.adder.in0[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B (.DIODE(\dpath.alu.adder.in1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__A (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__B (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__B (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__A (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__B (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B (.DIODE(\dpath.alu.adder.in1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A (.DIODE(\dpath.alu.adder.in0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__B (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(\dpath.alu.adder.in0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__C (.DIODE(_01875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__D (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__C (.DIODE(_01940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__A (.DIODE(\ctrl.d2c_inst[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__B (.DIODE(\ctrl.d2c_inst[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__C (.DIODE(\ctrl.d2c_inst[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__D (.DIODE(\ctrl.d2c_inst[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B (.DIODE(\ctrl.d2c_inst[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A1 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__B2 (.DIODE(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A1 (.DIODE(\ctrl.d2c_inst[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A1 (.DIODE(\ctrl.d2c_inst[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__B (.DIODE(net3436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B (.DIODE(net3307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B (.DIODE(net3424));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__B (.DIODE(net3312));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A (.DIODE(net3202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A (.DIODE(net3392));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(net3452));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A (.DIODE(net3420));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A (.DIODE(net3421));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A (.DIODE(net3461));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__A (.DIODE(net3435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__A (.DIODE(net3216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__07471__B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__B (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__B (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__S (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07502__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__S (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07515__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__S (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__S (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__B (.DIODE(net3308));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A0 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__S (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__S (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__S (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__S (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__S (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A1 (.DIODE(\dpath.RF.wdata[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__S (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__S (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07695__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__S (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__S (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07734__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__S (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__S (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__S (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__S (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__S (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__S (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__S (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__C1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__B1 (.DIODE(_01804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A1 (.DIODE(\ctrl.d2c_inst[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__B2 (.DIODE(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__B1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A (.DIODE(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__B2 (.DIODE(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A1 (.DIODE(\ctrl.d2c_inst[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A1 (.DIODE(\ctrl.d2c_inst[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__B (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A2 (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__B (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__B (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__C (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__D (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A2 (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B2 (.DIODE(_02099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A1 (.DIODE(net3202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__B (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B2 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__B1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__C1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A2 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__B (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__C (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__D (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__C (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__D (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A1_N (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A2_N (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__S (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A2 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__B (.DIODE(net3273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__B (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__B1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__C1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__B (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__C (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__B1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__B2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__B (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__B (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__B1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A2 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__B (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__B (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__C (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__B1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__B1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B2 (.DIODE(_02284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__C (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A2 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__A (.DIODE(net3392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A (.DIODE(net3392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A2 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__C1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__S0 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__S1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B2 (.DIODE(_02347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__B1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__B2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__C (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__D (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__C (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__B1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__B2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__C1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A (.DIODE(net3452));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__A (.DIODE(net3452));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__B (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__C1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__D (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__A1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B2 (.DIODE(_01785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__B (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__A (.DIODE(net3420));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__A (.DIODE(net3420));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__B1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__C1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__S0 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__B1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__B (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__C (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__B2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__C (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__D (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__B (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A2 (.DIODE(_02551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08344__A (.DIODE(net3421));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A (.DIODE(net3421));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A2 (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A2 (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B1 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__C1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__B2 (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__C (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__D (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__B (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__C (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__B2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__B2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A (.DIODE(net3461));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A (.DIODE(net3461));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A2 (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A2 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__B (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__C1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__S0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__S1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__B1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__B2 (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__B1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__B2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__A1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__C (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__D (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A2 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__B2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__C1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__B (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net3435));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A (.DIODE(net3435));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A2 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__S0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__S1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__B1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__B2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__B (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__C (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__B1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__C (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__D (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__B2 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__B (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__C1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A2 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__B1_N (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08643__A2_N (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08643__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__A2 (.DIODE(_02841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__B1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__B2 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__B1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__D (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__B2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__B (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__D (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__A1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__B2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__C (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__B (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A2 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__B (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A2 (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__B (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__C (.DIODE(_02947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__A2_N (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A2 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__S0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__S1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__08764__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__B1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__B1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__B2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__B (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__C (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A1 (.DIODE(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__B2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__B (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__B (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__C (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__D (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__A1 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__B1 (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__B (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__D (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A1 (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__B (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__C1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__A2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__B1 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A2 (.DIODE(_03054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__C (.DIODE(_03054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__B1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08860__A1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08860__A2 (.DIODE(_03053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__S0 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__S1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__B1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__08880__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__B2 (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__B (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__B1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__C (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__B2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__B (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__A (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__C (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__D (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__B (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__B (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__B2 (.DIODE(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__B2 (.DIODE(net765));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__C (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__D (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__B (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__C1 (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A2 (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__B (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__A2_N (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A2 (.DIODE(_03167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A1 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__C1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__S0 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__S1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A1 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__B1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A1 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__C1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__B1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__B2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__B (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09002__B (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__B1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__C (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__B (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__C (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__D (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A2 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__B1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__D (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09044__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09044__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A1_N (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__B1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A2 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__C1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__B2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__B1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__C (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__B1 (.DIODE(\dpath.alu.adder.in0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__B2 (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__C (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__D (.DIODE(\dpath.alu.adder.in0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__B (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__A (.DIODE(net788));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__B (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__B2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__C (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__D (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__A (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__B1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__A1 (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A (.DIODE(_03410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__B1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A2 (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__C1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__S0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__S1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__B1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__B2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__B (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__C (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__B2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__D (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__C (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__D (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__B (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A2 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__B2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__C (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__D (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__A1 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__B (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__C1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A1 (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__B1 (.DIODE(_03446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__B (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__B1 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A2 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__C1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A2 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__B (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__B (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__C (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__D (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__B2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A2 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B1 (.DIODE(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__C (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__D (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B1 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A2 (.DIODE(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__B (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__C (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__B2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__D (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A1 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__B1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__B1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A2 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__C1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__B2 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__B (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__C (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__D (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__B2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A2 (.DIODE(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__C (.DIODE(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__D (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__B (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A2 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__B2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A1 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__D (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__D (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__C1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A1 (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A2 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B1 (.DIODE(_02946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A2 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B2 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__C1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__B (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A2 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__C (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__D (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A1 (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__A2 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__B2 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__B1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__C (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__D (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__B (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__B (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A2 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__B2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__A (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__D (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__C (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A1_N (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A2_N (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A2 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__B (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__C (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__D (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B2 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__B2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__C (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__D (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A2 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__B (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__A (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A1 (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A2 (.DIODE(_03968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A2 (.DIODE(_03969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09792__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__C1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__S0 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__S1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A2 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__C (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__D (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A1_N (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A2_N (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__D (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__C (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__D (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A1 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A2 (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__B2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__B (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__C (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A2 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__B2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__D (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A2 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__B (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__C (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__B2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A3 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A4 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A2 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__B1 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__B (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__C (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__D (.DIODE(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__A1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__B1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__C1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A1 (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A2 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__B (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__B1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__C1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__B1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__B2 (.DIODE(_04151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A2 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__B1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__C (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__D (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A1_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A2_N (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__D (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A (.DIODE(\dpath.alu.adder.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A1 (.DIODE(\dpath.alu.adder.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__A (.DIODE(\dpath.alu.adder.in1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A1 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A2 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A3 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A4 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__A1 (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__B2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A1 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A2 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__B (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__C (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__D (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__B1 (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__B2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__D (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A1_N (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A2_N (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__C (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__D (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__A1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__A2 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__B2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__D (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__A (.DIODE(\dpath.alu.adder.in0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__B (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__D (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__B (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__B1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__B2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__C (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__D (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__B (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__B2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__A2 (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__B1 (.DIODE(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__B2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__B1 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A2 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A2 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__B (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__S0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__S1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__C1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__B1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__B2 (.DIODE(_04301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__D (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__B1 (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__B2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__B (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__A1 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__A2 (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__C (.DIODE(\dpath.alu.adder.in1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__D (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__A2 (.DIODE(\dpath.alu.adder.in1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__B1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__B2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__B (.DIODE(\dpath.alu.adder.in1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__A1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__C (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A1 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B2 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__B (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__B (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__C (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A2 (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__B1 (.DIODE(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__B2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A (.DIODE(_04335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__B1 (.DIODE(_04335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__B2 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__C (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__D (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A1_N (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A2_N (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__A (.DIODE(\dpath.alu.adder.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A2 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__B (.DIODE(\dpath.alu.adder.in0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__A (.DIODE(\dpath.alu.adder.in1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__B (.DIODE(\dpath.alu.adder.in0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__C (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__D (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__B2 (.DIODE(net766));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A1 (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__B1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__A2 (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A2 (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__B1 (.DIODE(_04302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A1 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__C1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__A (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__A (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__A1 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__B1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__10257__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__B2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A2 (.DIODE(\dpath.alu.adder.in1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__B1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__B2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__C (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A (.DIODE(\dpath.alu.adder.in1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__B (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__B1 (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__B2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__B (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__C (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__D (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A2 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__B2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__C (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__C (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__D (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__A1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__A2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__C (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__D (.DIODE(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A2 (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__B1 (.DIODE(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__B2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__B (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__C (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A1 (.DIODE(net773));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__B1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__B2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__B (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A2 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A3 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A4 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A1 (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A2 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__C (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__D (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A2 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__B2 (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__A (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__B1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A2 (.DIODE(_04593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__B1 (.DIODE(_04453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__B (.DIODE(net3542));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B (.DIODE(net3542));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__B1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A2 (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A1 (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A1 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__C1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__S0 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__S1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__S0 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__S1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__A1 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A (.DIODE(_02097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__B2 (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A2 (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__B1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__B2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__B2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__C (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__B2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__C (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A2 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__B (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__C (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__D (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__B (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__C (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__D (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__B1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__B2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__B (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__B (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__B1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__B2 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__C_N (.DIODE(_04675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B1_N (.DIODE(_04675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__C (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__D (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__B2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A1 (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A2 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__B (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A2 (.DIODE(\dpath.alu.adder.in0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__B (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__B (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A2 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__B2 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__C (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__D (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__B1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__B2 (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__C1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A2 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A2 (.DIODE(_04760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__C1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__B1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__B2 (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__B (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__B1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__B2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__C (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__D (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A1_N (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A2_N (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__C (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__D (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__B2 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__B2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__C (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__D (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__B2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__C (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__D (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__C (.DIODE(\dpath.alu.adder.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__D (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__C (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__D (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A1 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A2 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__B1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__B2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A2 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__B2 (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__B1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__B2 (.DIODE(\dpath.alu.adder.in0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B1 (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__C (.DIODE(\dpath.alu.adder.in0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__D (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__A2 (.DIODE(\dpath.alu.adder.in0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__B2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__B (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__B (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__B (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__B (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__B2 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__C (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__D (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A2 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__B1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__B2 (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A1 (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__B1 (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__A2 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10743__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A2 (.DIODE(net3542));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A2 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10756__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__C1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__B1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__B2 (.DIODE(_04968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A2 (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__B1 (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__B2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__B (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__C (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__B1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__B2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__C (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A1 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__A1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__C (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__D (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__C (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__D (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__B2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__C (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__B (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__C (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__D (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A (.DIODE(\dpath.alu.adder.in1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__C (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__D (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A1 (.DIODE(\dpath.alu.adder.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A2 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__B2 (.DIODE(\dpath.alu.adder.in1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__B (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A2 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10840__B (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A2 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B1 (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__B (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__C (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__D (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A1 (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__B1 (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__B2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__B (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__B (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__B (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__C (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__D (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__B2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A2 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__S (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__B1 (.DIODE(_01875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__A1 (.DIODE(_01875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A2 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__B (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__S0 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__S1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__C1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__S (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B2 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A (.DIODE(_01875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A2 (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B1 (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A1 (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__B (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__B2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__B1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__B2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__C (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__D (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__B2 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__C (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__B2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__B1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__C (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__A1 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__A1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__A2 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__B2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__C (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__D (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__C (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__D (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__B (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__B1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__B2 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__C (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__D (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A2 (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B1 (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__B (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A2 (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__B (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__B (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__B (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A1 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A2 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A3 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A4 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A2 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__B2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__B2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__C (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__D (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__C1 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A1 (.DIODE(_01787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__B (.DIODE(_05293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__B1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__C1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__B1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__B2 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B (.DIODE(\dpath.alu.adder.in1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A2 (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__B1 (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__B2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__C (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__D (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__B (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__A1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__A2 (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__B2 (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__B1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__B2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__C (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__D (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__C (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__B2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A2 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__C (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A2 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__B2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__C (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__D (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A1 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__A1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__A2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__B1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__A2 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A2 (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B1 (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__C (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__D (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A1_N (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A2_N (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__C (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__D (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__B (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B (.DIODE(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__B (.DIODE(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__B2 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A2 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__B2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__C (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__D (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A2 (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__B (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A0 (.DIODE(net3674));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__S (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__S (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A1 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__B (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__B (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__C1 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11302__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__11302__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__B1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__S0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__S1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__C1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11314__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11314__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__S0 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__S1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__B1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A2 (.DIODE(_02115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B1 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B2 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A1 (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A2 (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__B1 (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__B2 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__C (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__D (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__B (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__B (.DIODE(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B (.DIODE(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__B2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A1 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__B1 (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__B2 (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__C (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__D (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__B (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A2 (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A1 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B2 (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__B (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__C (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__D (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A2 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B2 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__B (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__C (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__D (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__B (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__B1 (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__B (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__C (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__D (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A2 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__A1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__A2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__B1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__B2 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__C (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__D (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__B1 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__B2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__C (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__D (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A1 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A2 (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B1 (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__B (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__C (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__D (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__A1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__A2 (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__B (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__B (.DIODE(\dpath.alu.adder.in1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__B (.DIODE(\dpath.alu.adder.in1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__B1 (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__B2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__C (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__D (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A2 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A (.DIODE(_02239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A1 (.DIODE(net3336));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__B (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__C1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__B1 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__B1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__B1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__S0 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__S1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__S0 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__S1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__C1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__A1 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A1 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__C1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A2 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__B2 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B (.DIODE(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__A (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__B (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__B1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__C1 (.DIODE(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A2 (.DIODE(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__A (.DIODE(net764));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B (.DIODE(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__B (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A2 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__B1 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__C1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__B (.DIODE(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A1 (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A2 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A1 (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A2 (.DIODE(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__A1 (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__B (.DIODE(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__A (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__B (.DIODE(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__B (.DIODE(\dpath.alu.adder.in0[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__B (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__B (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__B (.DIODE(\dpath.alu.adder.in1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__B (.DIODE(\dpath.alu.adder.in1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__B (.DIODE(\dpath.alu.adder.in1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A2 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__B (.DIODE(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__B (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__B (.DIODE(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__B (.DIODE(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__B (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__11614__A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA__11614__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A1 (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A2 (.DIODE(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A2 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__C1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A2 (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A1 (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A2 (.DIODE(_05828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__B (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__B1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__B2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__C1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__S (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11681__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__S (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11687__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__11697__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11699__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__S (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11723__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(\dpath.RF.wdata[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__S (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A0 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11737__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__S (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A0 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__A0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11761__S (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__S (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__S (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11806__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__S (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11816__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__A1 (.DIODE(\dpath.RF.wdata[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__S (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__S (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__S (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11872__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__S (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__S (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__S (.DIODE(_05851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__A0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__S (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__A0 (.DIODE(\dpath.RF.wdata[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__S (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__11929__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A0 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__S (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A0 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A0 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11948__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__A0 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A0 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11956__A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__11956__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A0 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__S (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11960__A0 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11960__S (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11962__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11964__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11966__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__S (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11982__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11986__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(\dpath.RF.wdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11992__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__S (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A0 (.DIODE(net3214));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12001__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A0 (.DIODE(net3257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A0 (.DIODE(net3443));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A0 (.DIODE(net3481));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A0 (.DIODE(net3523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__A0 (.DIODE(net3516));
 sky130_fd_sc_hd__diode_2 ANTENNA__12011__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__A0 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A0 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A0 (.DIODE(net3497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A0 (.DIODE(net3502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__A0 (.DIODE(net3512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__A0 (.DIODE(\dpath.csrw_out0.d[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12024__A0 (.DIODE(\dpath.csrw_out0.d[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__A0 (.DIODE(net3433));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__A0 (.DIODE(net3457));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__A0 (.DIODE(net3404));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__A0 (.DIODE(net3366));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__A0 (.DIODE(net3334));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__A0 (.DIODE(net3247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__A0 (.DIODE(net3488));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__A0 (.DIODE(net3486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12042__A0 (.DIODE(net3500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__A0 (.DIODE(net3448));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__A0 (.DIODE(net3255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A0 (.DIODE(net3217));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A0 (.DIODE(net3450));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A0 (.DIODE(net3430));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A0 (.DIODE(net3380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__A0 (.DIODE(net3459));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__S (.DIODE(_05860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__A0 (.DIODE(net3437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A0 (.DIODE(net3505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A0 (.DIODE(net3289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__S (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12066__A (.DIODE(net3214));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__A (.DIODE(net3257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__A (.DIODE(\dpath.csrw_out0.d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__A (.DIODE(\dpath.csrw_out0.d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__A (.DIODE(\dpath.csrw_out0.d[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__C (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A (.DIODE(\dpath.csrw_out0.d[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A (.DIODE(\dpath.csrw_out0.d[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A (.DIODE(\dpath.csrw_out0.d[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A (.DIODE(\dpath.csrw_out0.d[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A (.DIODE(\dpath.csrw_out0.d[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A (.DIODE(\dpath.csrw_out0.d[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__C1 (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__A (.DIODE(\dpath.csrw_out0.d[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A (.DIODE(net3247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__A (.DIODE(\dpath.csrw_out0.d[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12105__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__A (.DIODE(\dpath.csrw_out0.d[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A (.DIODE(\dpath.csrw_out0.d[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__A (.DIODE(\dpath.csrw_out0.d[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__A (.DIODE(net3255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12113__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__A (.DIODE(net3217));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__A (.DIODE(\dpath.csrw_out0.d[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A (.DIODE(\dpath.csrw_out0.d[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__C1 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A (.DIODE(net3380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__A (.DIODE(\dpath.csrw_out0.d[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__C1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__A (.DIODE(\dpath.csrw_out0.d[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__C1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__A (.DIODE(\dpath.csrw_out0.d[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__C1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A (.DIODE(net3289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__C (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__C1 (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A1 (.DIODE(net3214));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1 (.DIODE(net3257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A1 (.DIODE(net3443));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__A1 (.DIODE(net3481));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A1 (.DIODE(net3523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A1 (.DIODE(net3516));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__A1 (.DIODE(net3548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__A1 (.DIODE(net3529));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A1 (.DIODE(net3497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__A1 (.DIODE(net3502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__A1 (.DIODE(net3512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A1 (.DIODE(\dpath.csrw_out0.d[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__A1 (.DIODE(\dpath.csrw_out0.d[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A1 (.DIODE(net3433));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__A1 (.DIODE(net3457));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A1 (.DIODE(net3404));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__C1 (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__A1 (.DIODE(net3366));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A1 (.DIODE(net3334));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A1 (.DIODE(net3247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__A1 (.DIODE(net3488));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__A1 (.DIODE(net3486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A1 (.DIODE(net3500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__A1 (.DIODE(net3448));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__A1 (.DIODE(net3255));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A1 (.DIODE(net3217));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A1 (.DIODE(net3450));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A1 (.DIODE(net3430));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__A1 (.DIODE(net3380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A1 (.DIODE(net3459));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A1 (.DIODE(net3437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A1 (.DIODE(net3505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A1 (.DIODE(net3289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__S (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__B1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__C1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__S (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__S (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__B1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__C1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__S1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__S0 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A_N (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B_N (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A0 (.DIODE(net3652));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__S (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__B (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__B1 (.DIODE(_05989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__B2 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__B (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__S (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__S (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__S (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__S (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__B1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__C1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__S0 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__S1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__S0 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__S1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A1 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__B1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__B2 (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__S (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A1 (.DIODE(net786));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B1 (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__B1 (.DIODE(net3682));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__B2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__S (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__A2 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__B1 (.DIODE(_06022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__B2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__B (.DIODE(_06024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__B (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__B (.DIODE(net3273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__B (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__B (.DIODE(net3400));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__B (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__B (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__B (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__B (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__B (.DIODE(_03053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__B (.DIODE(_03167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__B (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__B (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__B (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__B (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__B (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__B (.DIODE(_03969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__B (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__B (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__B (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__B (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__B (.DIODE(_04760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__B (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__B (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__B (.DIODE(_05293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__B (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__B (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__B (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A2 (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A_N (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__C (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__S0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__S0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__S1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__B1_N (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__B (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A1 (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__C1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__A1 (.DIODE(_05989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__A1 (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__S0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__C1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__B1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12350__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__S (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__B (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__C (.DIODE(_06022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A1 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__B1 (.DIODE(_06089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__S0 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__S1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__S0 (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__S1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__C1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__S0 (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__S1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__S (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12373__S (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__B1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__S (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__B (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__C (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A1 (.DIODE(_02099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A2 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__A1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__C1 (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__S (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__S (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__B1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__S (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__S (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A1 (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A1_N (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__B1 (.DIODE(_06135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__S (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__S (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__B1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12415__S (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__S (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__B2 (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A1 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__A1_N (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__B1 (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__S (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__S (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__B1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__S (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__B2 (.DIODE(_02284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A1 (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__A1_N (.DIODE(net3392));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__B1 (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__S (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__S (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__B1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__S (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__S0 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__S1 (.DIODE(net801));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__B2 (.DIODE(_02347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__A1_N (.DIODE(net3452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__B1 (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__S (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__S (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__B1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__S (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__S (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__S0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A1_N (.DIODE(net3420));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B1 (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12510__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__B1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12516__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__B1 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__C1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__C_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__S0 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__S0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__S1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A1 (.DIODE(_02551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12530__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A1_N (.DIODE(net3421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__B1 (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__B1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__S (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__S (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__B1 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__A1 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__C1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__C_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__S0 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__S1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B2 (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__A1 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A1_N (.DIODE(net3461));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__B1 (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__S (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__B1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__S (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__B1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__C1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__C_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__S0 (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__S1 (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__S0 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__S1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__B2 (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A1_N (.DIODE(net3435));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A2_N (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__S (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__S (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__B1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__S (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__S (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__C1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__S0 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__S1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__S0 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__A1 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A2 (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__B1 (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12608__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12608__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__S (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__B1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__S0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__B2 (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A2 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__S (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__S (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__B1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__A1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__S (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__S (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A1 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__B1 (.DIODE(net796));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__C1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__C_N (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__S0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12651__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A1 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__A2 (.DIODE(_06375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__S (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__S (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__S0 (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__S1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__S (.DIODE(net826));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__S (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__B1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__C1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__C_N (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__S0 (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__S0 (.DIODE(net823));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__S1 (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__S0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__S1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__B2 (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A1 (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A2 (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12682__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__B1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__A1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__C1 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__S1 (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__B1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__C1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__S0 (.DIODE(net822));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__S1 (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__S0 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__S1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__A2 (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__S0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A2 (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__S (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__S (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__S0 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__S1 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__S0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A2 (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__S (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__S (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12775__S0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12775__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12777__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A2 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12783__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__S (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__S0 (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__S0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__B2 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A2 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__S (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__S0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A1 (.DIODE(_03968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A2 (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__S (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__S (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__S (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__S0 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__S1 (.DIODE(net811));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__S0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A1 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__A2 (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__B1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12865__S (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__S (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__A1 (.DIODE(_01788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__B1 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__A1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__C1 (.DIODE(_01790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12870__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__S0 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12877__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__B2 (.DIODE(_04151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__A1 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__A2 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__B1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__B1 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__C_N (.DIODE(net3665));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__S0 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__S1 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__S0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__B2 (.DIODE(_04301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A1 (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A2 (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__S (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__S (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__B1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12913__A1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12913__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12915__S (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__S (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__B1 (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__C_N (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__S0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__S1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__B2 (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A1 (.DIODE(_04593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A2 (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__B1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__S1 (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__S (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__C1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__12945__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12947__S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__S0 (.DIODE(net834));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__S0 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__S1 (.DIODE(net812));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__S0 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__B2 (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A2 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A2 (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__B1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__S0 (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__S0 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__B2 (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A1 (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B1 (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__B1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__C1 (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A1 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__S0 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__B2 (.DIODE(_04968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A1 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__B1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__C1 (.DIODE(net3669));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__S0 (.DIODE(net838));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__S1 (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__S0 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__A2 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__B2 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__A1 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A1 (.DIODE(_01975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__B1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__B1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__C1 (.DIODE(net3669));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__S (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__S (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__S0 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__B2 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A1 (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__A1 (.DIODE(_01975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__B1 (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__B1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__C1 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__S (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__C_N (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__S0 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__S0 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__S1 (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__S0 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13076__A (.DIODE(net3665));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__B2 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__A1 (.DIODE(_05662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__B1 (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__S (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__S (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__B1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__A1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__A1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__C1 (.DIODE(net3669));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__S0 (.DIODE(net840));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__S (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__S (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__A1 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__B1 (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A1 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__C1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__C_N (.DIODE(net3665));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__S1 (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__S0 (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__S1 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__S0 (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__S1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B1 (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B2 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A1 (.DIODE(_05828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__B1 (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13138__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13139__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__B (.DIODE(_06089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__B (.DIODE(_06135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__B (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__B (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__B (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__B (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__B (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__B (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__B (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__B (.DIODE(_06375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__B (.DIODE(_06399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__B (.DIODE(_06423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__B (.DIODE(_06447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__B (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__B (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__B (.DIODE(_06543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__B (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__B (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__B (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__B (.DIODE(_05989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__B (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__B (.DIODE(_02099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__B (.DIODE(_02217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B (.DIODE(_02284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__B (.DIODE(_02347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__B (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__B (.DIODE(_02874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__B (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__B (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__B (.DIODE(_04151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__B (.DIODE(_04301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__B (.DIODE(_04452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13197__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13197__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__B (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__B (.DIODE(_04968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__B (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__B (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__B (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__B (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13211__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13220__S (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13224__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13228__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__A1 (.DIODE(\dpath.RF.wdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__S (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__A (.DIODE(\ctrl.d2c_inst[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__A (.DIODE(\ctrl.d2c_inst[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__B (.DIODE(\ctrl.d2c_inst[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__C (.DIODE(\ctrl.d2c_inst[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__D (.DIODE(\ctrl.d2c_inst[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__A (.DIODE(\ctrl.d2c_inst[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__B (.DIODE(\ctrl.d2c_inst[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__13245__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__13247__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__13248__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13249__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__13250__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__13251__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__13257__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__13263__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13276__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__13278__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13282__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__13284__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13285__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__13287__A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__B1 (.DIODE(_06846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13290__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__13292__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__13295__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13297__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__13298__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__13299__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__13301__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13303__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__13304__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13306__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__13307__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13309__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__13313__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13315__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__13317__A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13327__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__13331__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__A2 (.DIODE(_06813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__B1 (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13343__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13357__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA__13361__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13366__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13369__A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__13371__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__13373__A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__13374__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13374__B (.DIODE(_05987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13375__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13375__B (.DIODE(_06022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__B (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__B (.DIODE(_02183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__B (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__B (.DIODE(_02316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__B (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13381__A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA__13381__B (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__B (.DIODE(_02551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13383__B (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__B (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__B (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__B (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__B (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__B (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__B (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__B (.DIODE(_03410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__B (.DIODE(net3673));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__B (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__A (.DIODE(net848));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__B (.DIODE(_03968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__B (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__B (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__B (.DIODE(_04593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__B (.DIODE(net3692));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__B (.DIODE(net3647));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__A1 (.DIODE(_06024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__S (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13410__A1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13410__S (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13411__A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__B (.DIODE(net3273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13414__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13416__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13416__B (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__B (.DIODE(net3400));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13423__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__B (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__B (.DIODE(_02841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__B (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A1 (.DIODE(_03053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__B (.DIODE(_03167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A1 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__B (.DIODE(net3454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A1 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__B (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__B (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__B (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13446__B (.DIODE(_03969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__B (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__B (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13451__A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__B (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13453__A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__A0 (.DIODE(net3542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__A1 (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__S (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13455__A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__B (.DIODE(_04760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A1 (.DIODE(_04934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__S (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__B (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__A1 (.DIODE(_05293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__S (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__B (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__B (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__A2 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__B (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13470__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__13478__A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__13479__A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA__13503__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__A0 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13505__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13507__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13508__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13509__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13513__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13514__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13517__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13518__S (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__13519__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13527__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__A0 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__A0 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__A0 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13533__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__A0 (.DIODE(\dpath.RF.wdata[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__S (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13538__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__13538__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13540__A0 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13540__S (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__C1 (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA__13550__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13551__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__13556__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__13556__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13565__C1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13569__A2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__B (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13574__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13585__A1 (.DIODE(net3542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__B (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A2 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__C1 (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13614__C1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA__13615__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__A1 (.DIODE(net3202));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13618__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__C1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13622__C1 (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13630__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__13630__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__B (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__A1 (.DIODE(net3392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13638__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__13639__A1 (.DIODE(net3452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13639__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__A1 (.DIODE(net3420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13642__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__A1 (.DIODE(net3421));
 sky130_fd_sc_hd__diode_2 ANTENNA__13643__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13644__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__A1 (.DIODE(net3461));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__A1 (.DIODE(net3435));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__A1 (.DIODE(net3216));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__C1 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA__13651__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__A1 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13653__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13654__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13655__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13657__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13659__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13661__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13663__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__S (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13667__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13668__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13669__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13672__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13674__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13676__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__13676__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13678__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__A1 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13682__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__13682__S (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13684__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13685__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13688__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13690__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__A1 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13693__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13695__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13696__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__S (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13700__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13702__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__13702__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13703__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__A1 (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__S (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__13715__A1 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__13715__S (.DIODE(_01742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13718__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13719__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13725__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13727__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13728__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13729__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13730__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13731__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__A1 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__S (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__A1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13736__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13737__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13739__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13740__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__A1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13743__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__A1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__S (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__B (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__13751__A2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__13752__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__A2_N (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__B1 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__A1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__A2 (.DIODE(_06024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13788__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13790__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13791__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__A2 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA__14581__CLK (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__14909__D (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14910__D (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14917__D (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14919__D (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14921__D (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14923__D (.DIODE(_01135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14925__D (.DIODE(_01137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14927__D (.DIODE(_01139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__D (.DIODE(_01140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__D (.DIODE(_01141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__D (.DIODE(_01142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14931__D (.DIODE(_01143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14932__D (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14933__D (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14934__D (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14935__D (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__D (.DIODE(_01148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14937__D (.DIODE(_01149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14939__D (.DIODE(_01151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15005__D (.DIODE(_01217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15007__D (.DIODE(_01219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15013__D (.DIODE(_01225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__D (.DIODE(_01242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15189__D (.DIODE(_01401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15190__D (.DIODE(_01402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15207__D (.DIODE(_01419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15209__D (.DIODE(_01421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__D (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__D (.DIODE(_01423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15215__D (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15216__D (.DIODE(_01428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15217__D (.DIODE(_01429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15218__D (.DIODE(_01430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15219__D (.DIODE(_01431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__D (.DIODE(_01432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15231__D (.DIODE(net3171));
 sky130_fd_sc_hd__diode_2 ANTENNA__15232__D (.DIODE(net3195));
 sky130_fd_sc_hd__diode_2 ANTENNA__15233__D (.DIODE(_01445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__D (.DIODE(net2093));
 sky130_fd_sc_hd__diode_2 ANTENNA__15235__D (.DIODE(_01447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15236__D (.DIODE(net3179));
 sky130_fd_sc_hd__diode_2 ANTENNA__15238__D (.DIODE(_01450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15240__D (.DIODE(net1971));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0__f_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10__f_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11__f_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12__f_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13__f_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14__f_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15__f_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1__f_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2__f_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3__f_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4__f_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5__f_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6__f_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7__f_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8__f_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9__f_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_A (.DIODE(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_A (.DIODE(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_clk_A (.DIODE(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_clk_A (.DIODE(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(_06063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(_02115_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(_02097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(_01685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(_02025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(_02025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(_02021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout396_A (.DIODE(_02021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout397_A (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout399_A (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(_01952_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(_01834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(_01833_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(_01833_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_A (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(_01822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(_01822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(_01743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(_01743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(_01742_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(_01741_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(_01741_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(_05851_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(_05849_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(_05849_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(_02026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout444_A (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout445_A (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_A (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout449_A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout450_A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout452_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(_01824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout456_A (.DIODE(_01824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(_05860_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(_01825_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(_01825_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(_02100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(_02100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(_02844_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout477_A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(_01975_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(_01804_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_A (.DIODE(_01804_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout482_A (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout483_A (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_A (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout489_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout491_A (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout492_A (.DIODE(_01790_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout493_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_A (.DIODE(_01790_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout495_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout496_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout498_A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout499_A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout500_A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout501_A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout502_A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout503_A (.DIODE(_01788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(_01788_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout506_A (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout507_A (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout508_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout509_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout510_A (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout511_A (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout512_A (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout513_A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout514_A (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout515_A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout516_A (.DIODE(_01771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout517_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout518_A (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout519_A (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_A (.DIODE(_00009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout523_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout524_A (.DIODE(_00008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout525_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout526_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout527_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout528_A (.DIODE(_00008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout529_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout530_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout532_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout533_A (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout534_A (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout535_A (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout536_A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout539_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout540_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout541_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout542_A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout543_A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout544_A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout545_A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout547_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout548_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout549_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout550_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout551_A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout552_A (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout553_A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout554_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout555_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout556_A (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout557_A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout558_A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout559_A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout560_A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout562_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout563_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout564_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout565_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout566_A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout567_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout568_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout569_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout570_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout571_A (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout572_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout573_A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout575_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout576_A (.DIODE(_00005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout577_A (.DIODE(net3216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout578_A (.DIODE(net3216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout579_A (.DIODE(\dpath.alu.adder.in0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout580_A (.DIODE(\dpath.alu.adder.in0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout581_A (.DIODE(\dpath.alu.adder.in0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout582_A (.DIODE(\dpath.alu.adder.in0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout583_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout585_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout590_A (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout592_A (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout593_A (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(\dpath.alu.adder.in0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout595_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout598_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(_06813_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout602_A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(\dpath.alu.adder.in0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(\dpath.alu.adder.in0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(\dpath.alu.adder.in0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(\dpath.alu.adder.in0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout613_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout614_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_A (.DIODE(\dpath.alu.adder.in0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(\dpath.alu.adder.in0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(\dpath.alu.adder.in0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_A (.DIODE(\dpath.alu.adder.in0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(\dpath.alu.adder.in0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout625_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout627_A (.DIODE(\dpath.alu.adder.in0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_A (.DIODE(\dpath.alu.adder.in0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_A (.DIODE(\dpath.alu.adder.in0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout630_A (.DIODE(\dpath.alu.adder.in0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout631_A (.DIODE(\dpath.alu.adder.in0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout632_A (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout633_A (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout634_A (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout635_A (.DIODE(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout636_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout637_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout638_A (.DIODE(\dpath.alu.adder.in0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout639_A (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout640_A (.DIODE(\dpath.alu.adder.in0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout641_A (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout642_A (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout643_A (.DIODE(\dpath.alu.adder.in0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout644_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout645_A (.DIODE(\dpath.alu.adder.in0[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout646_A (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout647_A (.DIODE(\dpath.alu.adder.in0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout648_A (.DIODE(\dpath.alu.adder.in0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout649_A (.DIODE(\dpath.alu.adder.in0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout650_A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout651_A (.DIODE(\dpath.alu.adder.in0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout652_A (.DIODE(\dpath.alu.adder.in0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout653_A (.DIODE(\dpath.alu.adder.in0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout654_A (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout655_A (.DIODE(\dpath.RF.wdata[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout658_A (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout662_A (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout666_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout667_A (.DIODE(\dpath.RF.wdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout668_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout669_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout675_A (.DIODE(net676));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout682_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout688_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_A (.DIODE(_06813_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout704_A (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout712_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout716_A (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout720_A (.DIODE(\dpath.alu.adder.in1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout721_A (.DIODE(\dpath.alu.adder.in1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout722_A (.DIODE(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout723_A (.DIODE(\dpath.alu.adder.in1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout724_A (.DIODE(\dpath.alu.adder.in1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout725_A (.DIODE(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout726_A (.DIODE(\dpath.alu.adder.in1[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout727_A (.DIODE(\dpath.alu.adder.in1[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout728_A (.DIODE(net729));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout729_A (.DIODE(\dpath.alu.adder.in1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout730_A (.DIODE(\dpath.alu.adder.in1[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout731_A (.DIODE(\dpath.alu.adder.in1[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout732_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout733_A (.DIODE(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout734_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout735_A (.DIODE(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout736_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout737_A (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout739_A (.DIODE(\dpath.alu.adder.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout742_A (.DIODE(\dpath.alu.adder.in1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout743_A (.DIODE(\dpath.alu.adder.in1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout746_A (.DIODE(\dpath.alu.adder.in1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout752_A (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout754_A (.DIODE(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout755_A (.DIODE(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout756_A (.DIODE(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout758_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout760_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout761_A (.DIODE(net762));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout762_A (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout764_A (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout765_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout766_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout767_A (.DIODE(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout768_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout769_A (.DIODE(net770));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout770_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout772_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout773_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout774_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout776_A (.DIODE(\dpath.alu.adder.in1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout777_A (.DIODE(\dpath.alu.adder.in1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout778_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout779_A (.DIODE(\dpath.alu.adder.in1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout780_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout781_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout783_A (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout784_A (.DIODE(\dpath.alu.adder.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout785_A (.DIODE(\dpath.alu.adder.in1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout786_A (.DIODE(\dpath.alu.adder.in1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout787_A (.DIODE(\dpath.alu.adder.in1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout788_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout789_A (.DIODE(\dpath.alu.adder.in1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout790_A (.DIODE(net791));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout791_A (.DIODE(net3665));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout792_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout794_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout795_A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout796_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout797_A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout798_A (.DIODE(net799));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout799_A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout800_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout801_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout802_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout803_A (.DIODE(net804));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout804_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout805_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout806_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout807_A (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout808_A (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout809_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout810_A (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout811_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout812_A (.DIODE(net813));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout813_A (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout814_A (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout815_A (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout816_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout817_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout818_A (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout819_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout820_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout821_A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout822_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout823_A (.DIODE(net824));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout824_A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout825_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout826_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout827_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout828_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout829_A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout830_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout831_A (.DIODE(net832));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout832_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout833_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout834_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout835_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout836_A (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout837_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout838_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout839_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout840_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout841_A (.DIODE(net842));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout842_A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout844_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout845_A (.DIODE(net846));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout846_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout847_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout848_A (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout849_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout850_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout851_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout852_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout853_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout855_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout857_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout858_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout859_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout860_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout861_A (.DIODE(net862));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout862_A (.DIODE(_01792_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout863_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout864_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout865_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout868_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout870_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout871_A (.DIODE(net872));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout872_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout873_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout874_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout875_A (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout876_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout877_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout878_A (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout879_A (.DIODE(_01792_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout880_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout881_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout882_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout883_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout884_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout886_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout887_A (.DIODE(net888));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout888_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout889_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout890_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout891_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout892_A (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout893_A (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout894_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1076_A (.DIODE(_01452_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1198_A (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2276_A (.DIODE(_01443_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2284_A (.DIODE(_01448_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2300_A (.DIODE(_01444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2331_A (.DIODE(\ctrl.d2c_inst[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2349_A (.DIODE(\dpath.sd_DX.q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2375_A (.DIODE(\dpath.sd_DX.q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2385_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2410_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2412_A (.DIODE(\ctrl.inst_X[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2413_A (.DIODE(\dpath.sd_DX.q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2416_A (.DIODE(_05991_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2417_A (.DIODE(\ctrl.inst_X[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2439_A (.DIODE(\dpath.csrw_out0.d[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2441_A (.DIODE(\dpath.csrr[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2442_A (.DIODE(_05662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2446_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2471_A (.DIODE(\dpath.csrw_out0.d[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2497_A (.DIODE(\ctrl.d2c_inst[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2505_A (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2509_A (.DIODE(\dpath.csrw_out0.d[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2520_A (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2522_A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2525_A (.DIODE(\ctrl.d2c_inst[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2526_A (.DIODE(\ctrl.d2c_inst[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2529_A (.DIODE(\ctrl.inst_X[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2535_A (.DIODE(\dpath.csrw_out0.d[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2538_A (.DIODE(\dpath.csrw_out0.d[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2540_A (.DIODE(\ctrl.d2c_inst[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2542_A (.DIODE(\dpath.csrw_out0.d[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2550_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2552_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2553_A (.DIODE(\dpath.csrw_out0.d[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2555_A (.DIODE(\dpath.csrw_out0.d[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2557_A (.DIODE(\ctrl.d2c_inst[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2559_A (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2562_A (.DIODE(\dpath.csrw_out0.d[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2564_A (.DIODE(\dpath.csrw_out0.d[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2566_A (.DIODE(\ctrl.d2c_inst[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2578_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2590_A (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2591_A (.DIODE(\dpath.csrw_out0.d[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2593_A (.DIODE(\dpath.csrw_out0.d[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2598_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2605_A (.DIODE(\dpath.csrw_out0.d[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2610_A (.DIODE(\dpath.csrw_out0.d[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2617_A (.DIODE(\dpath.csrw_out0.d[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2619_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2628_A (.DIODE(\dpath.csrw_out0.d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2632_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2646_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2653_A (.DIODE(\dpath.csrw_out0.d[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2674_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2678_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2692_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2694_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2695_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2696_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2701_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2703_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2707_A (.DIODE(_04933_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2710_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2711_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2715_A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2726_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2727_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2728_A (.DIODE(\dpath.RF.wdata[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2729_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2734_A (.DIODE(_02841_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2737_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2738_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2739_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2740_A (.DIODE(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2741_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2743_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2744_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2745_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2746_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2747_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2748_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2750_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2752_A (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2757_A (.DIODE(\dpath.csrr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2759_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2760_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2763_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2768_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2769_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2770_A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2772_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2774_A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2778_A (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2780_A (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2781_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2782_A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2785_A (.DIODE(_05828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2786_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2787_A (.DIODE(\dpath.csrr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2794_A (.DIODE(\dpath.RF.wdata[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2797_A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2850_A (.DIODE(\ctrl.d2c_inst[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2859_A (.DIODE(\ctrl.d2c_inst[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2861_A (.DIODE(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_output229_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_output239_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_output249_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_output250_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_output253_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_output254_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_output255_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_output256_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_output271_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_output330_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_output331_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_output332_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_output333_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_output347_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_output348_A (.DIODE(net348));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_203_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_204_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_208_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_211_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_211_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_997 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__conb_1 Proc_895 (.HI(net895));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06903_ (.A(net3349),
    .Y(_01749_));
 sky130_fd_sc_hd__inv_2 _06904_ (.A(net3285),
    .Y(_01750_));
 sky130_fd_sc_hd__inv_2 _06905_ (.A(net3403),
    .Y(_01751_));
 sky130_fd_sc_hd__inv_2 _06906_ (.A(net3393),
    .Y(_01752_));
 sky130_fd_sc_hd__inv_2 _06907_ (.A(net3432),
    .Y(_01753_));
 sky130_fd_sc_hd__inv_2 _06908_ (.A(\ctrl.d2c_inst[19] ),
    .Y(_01754_));
 sky130_fd_sc_hd__inv_2 _06909_ (.A(\ctrl.d2c_inst[18] ),
    .Y(_01755_));
 sky130_fd_sc_hd__inv_2 _06910_ (.A(\ctrl.d2c_inst[17] ),
    .Y(_01756_));
 sky130_fd_sc_hd__inv_2 _06911_ (.A(\ctrl.d2c_inst[16] ),
    .Y(_01757_));
 sky130_fd_sc_hd__inv_2 _06912_ (.A(\ctrl.d2c_inst[15] ),
    .Y(_01758_));
 sky130_fd_sc_hd__inv_2 _06913_ (.A(net3263),
    .Y(_01759_));
 sky130_fd_sc_hd__inv_2 _06914_ (.A(net3507),
    .Y(_01760_));
 sky130_fd_sc_hd__inv_2 _06915_ (.A(net242),
    .Y(_01761_));
 sky130_fd_sc_hd__inv_2 _06916_ (.A(net3325),
    .Y(_01762_));
 sky130_fd_sc_hd__inv_2 _06917_ (.A(net1156),
    .Y(_01763_));
 sky130_fd_sc_hd__inv_2 _06918_ (.A(net3309),
    .Y(_01764_));
 sky130_fd_sc_hd__inv_2 _06919_ (.A(net3243),
    .Y(_01765_));
 sky130_fd_sc_hd__inv_2 _06920_ (.A(net3245),
    .Y(_01766_));
 sky130_fd_sc_hd__inv_2 _06921_ (.A(net3281),
    .Y(_01767_));
 sky130_fd_sc_hd__inv_2 _06922_ (.A(net3279),
    .Y(_01768_));
 sky130_fd_sc_hd__inv_2 _06923_ (.A(net3259),
    .Y(_01769_));
 sky130_fd_sc_hd__inv_2 _06924_ (.A(net543),
    .Y(_01770_));
 sky130_fd_sc_hd__inv_4 _06925_ (.A(net535),
    .Y(_01771_));
 sky130_fd_sc_hd__inv_2 _06926_ (.A(net523),
    .Y(_01772_));
 sky130_fd_sc_hd__inv_2 _06927_ (.A(\ctrl.val_MW.q ),
    .Y(_01773_));
 sky130_fd_sc_hd__inv_2 _06928_ (.A(\ctrl.inst_W[3] ),
    .Y(_01774_));
 sky130_fd_sc_hd__inv_2 _06929_ (.A(\ctrl.inst_W[13] ),
    .Y(_01775_));
 sky130_fd_sc_hd__inv_2 _06930_ (.A(\ctrl.c2d_rf_waddr_W[0] ),
    .Y(_01776_));
 sky130_fd_sc_hd__inv_2 _06931_ (.A(\ctrl.c2d_rf_waddr_W[1] ),
    .Y(_01777_));
 sky130_fd_sc_hd__inv_2 _06932_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .Y(_01778_));
 sky130_fd_sc_hd__inv_2 _06933_ (.A(\ctrl.c2d_rf_waddr_W[3] ),
    .Y(_01779_));
 sky130_fd_sc_hd__inv_2 _06934_ (.A(\ctrl.c2d_rf_waddr_W[4] ),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_2 _06935_ (.A(net3203),
    .Y(_01781_));
 sky130_fd_sc_hd__inv_2 _06936_ (.A(net1172),
    .Y(_01782_));
 sky130_fd_sc_hd__inv_2 _06937_ (.A(net3200),
    .Y(_01783_));
 sky130_fd_sc_hd__inv_2 _06938_ (.A(net2950),
    .Y(_01784_));
 sky130_fd_sc_hd__inv_2 _06939_ (.A(net3399),
    .Y(_01785_));
 sky130_fd_sc_hd__inv_2 _06940_ (.A(net3631),
    .Y(_01786_));
 sky130_fd_sc_hd__inv_2 _06941_ (.A(net3609),
    .Y(_01787_));
 sky130_fd_sc_hd__inv_2 _06942_ (.A(net811),
    .Y(_01788_));
 sky130_fd_sc_hd__inv_6 _06943_ (.A(net799),
    .Y(_01789_));
 sky130_fd_sc_hd__inv_2 _06944_ (.A(net794),
    .Y(_01790_));
 sky130_fd_sc_hd__inv_2 _06945_ (.A(\ctrl.inst_W[20] ),
    .Y(_01791_));
 sky130_fd_sc_hd__clkinv_4 _06946_ (.A(net892),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(\ctrl.inst_M[1] ),
    .B(\ctrl.inst_M[0] ),
    .Y(_01793_));
 sky130_fd_sc_hd__or3_1 _06948_ (.A(\ctrl.inst_M[3] ),
    .B(\ctrl.inst_M[2] ),
    .C(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__or3b_1 _06949_ (.A(\ctrl.inst_M[12] ),
    .B(\ctrl.inst_M[14] ),
    .C_N(\ctrl.inst_M[13] ),
    .X(_01795_));
 sky130_fd_sc_hd__or3_1 _06950_ (.A(\ctrl.inst_M[6] ),
    .B(_01794_),
    .C(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__and3b_4 _06951_ (.A_N(_01796_),
    .B(_01769_),
    .C(\ctrl.inst_M[5] ),
    .X(net194));
 sky130_fd_sc_hd__and3_1 _06952_ (.A(\ctrl.inst_M[3] ),
    .B(\ctrl.inst_M[2] ),
    .C(\ctrl.inst_M[6] ),
    .X(_01797_));
 sky130_fd_sc_hd__or4bb_1 _06953_ (.A(_01793_),
    .B(\ctrl.inst_M[4] ),
    .C_N(\ctrl.inst_M[5] ),
    .D_N(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__nand2_1 _06954_ (.A(\ctrl.inst_M[5] ),
    .B(\ctrl.inst_M[6] ),
    .Y(_01799_));
 sky130_fd_sc_hd__or4_1 _06955_ (.A(\ctrl.inst_M[28] ),
    .B(\ctrl.inst_M[27] ),
    .C(\ctrl.inst_M[30] ),
    .D(\ctrl.inst_M[29] ),
    .X(_01800_));
 sky130_fd_sc_hd__o31a_1 _06956_ (.A1(\ctrl.inst_M[31] ),
    .A2(\ctrl.inst_M[26] ),
    .A3(_01800_),
    .B1(\ctrl.inst_M[5] ),
    .X(_01801_));
 sky130_fd_sc_hd__or4_1 _06957_ (.A(\ctrl.inst_M[6] ),
    .B(\ctrl.inst_M[12] ),
    .C(\ctrl.inst_M[13] ),
    .D(\ctrl.inst_M[14] ),
    .X(_01802_));
 sky130_fd_sc_hd__o22a_1 _06958_ (.A1(_01795_),
    .A2(_01799_),
    .B1(_01801_),
    .B2(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__o31a_4 _06959_ (.A1(_01769_),
    .A2(_01794_),
    .A3(_01803_),
    .B1(_01798_),
    .X(_01804_));
 sky130_fd_sc_hd__nor2_1 _06960_ (.A(\ctrl.inst_M[4] ),
    .B(\ctrl.inst_M[12] ),
    .Y(_01805_));
 sky130_fd_sc_hd__mux2_1 _06961_ (.A0(\ctrl.inst_M[12] ),
    .A1(_01805_),
    .S(\ctrl.inst_M[2] ),
    .X(_01806_));
 sky130_fd_sc_hd__or4b_1 _06962_ (.A(\ctrl.inst_M[13] ),
    .B(\ctrl.inst_M[14] ),
    .C(_01799_),
    .D_N(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__o31a_4 _06963_ (.A1(\ctrl.inst_M[3] ),
    .A2(_01793_),
    .A3(_01807_),
    .B1(_01804_),
    .X(net195));
 sky130_fd_sc_hd__or3_4 _06964_ (.A(_01778_),
    .B(\ctrl.c2d_rf_waddr_W[3] ),
    .C(\ctrl.c2d_rf_waddr_W[4] ),
    .X(_01808_));
 sky130_fd_sc_hd__nand2_1 _06965_ (.A(\ctrl.inst_W[1] ),
    .B(\ctrl.inst_W[0] ),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _06966_ (.A(\ctrl.inst_W[2] ),
    .B(\ctrl.inst_W[6] ),
    .Y(_01810_));
 sky130_fd_sc_hd__or4b_1 _06967_ (.A(\ctrl.inst_W[4] ),
    .B(_01809_),
    .C(_01810_),
    .D_N(\ctrl.inst_W[5] ),
    .X(_01811_));
 sky130_fd_sc_hd__or3_1 _06968_ (.A(\ctrl.inst_W[3] ),
    .B(\ctrl.inst_W[2] ),
    .C(_01809_),
    .X(_01812_));
 sky130_fd_sc_hd__nand3_1 _06969_ (.A(\ctrl.inst_W[5] ),
    .B(\ctrl.inst_W[6] ),
    .C(\ctrl.inst_W[12] ),
    .Y(_01813_));
 sky130_fd_sc_hd__or2_1 _06970_ (.A(_01812_),
    .B(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__or4b_1 _06971_ (.A(\ctrl.inst_W[4] ),
    .B(\ctrl.inst_W[6] ),
    .C(\ctrl.inst_W[12] ),
    .D_N(\ctrl.inst_W[5] ),
    .X(_01815_));
 sky130_fd_sc_hd__or4_1 _06972_ (.A(\ctrl.inst_W[14] ),
    .B(_01775_),
    .C(_01812_),
    .D(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__o31a_1 _06973_ (.A1(\ctrl.inst_W[3] ),
    .A2(\ctrl.inst_W[12] ),
    .A3(_01811_),
    .B1(_01814_),
    .X(_01817_));
 sky130_fd_sc_hd__o31ai_4 _06974_ (.A1(\ctrl.inst_W[14] ),
    .A2(\ctrl.inst_W[13] ),
    .A3(_01817_),
    .B1(_01816_),
    .Y(_01818_));
 sky130_fd_sc_hd__or2_2 _06975_ (.A(_01776_),
    .B(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__nor2_2 _06976_ (.A(_01777_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__or2_2 _06977_ (.A(_01777_),
    .B(_01819_),
    .X(_01821_));
 sky130_fd_sc_hd__or2_4 _06978_ (.A(_01808_),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _06979_ (.A0(net718),
    .A1(net2654),
    .S(net413),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _06980_ (.A0(net717),
    .A1(net3112),
    .S(net413),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _06981_ (.A0(net714),
    .A1(net3046),
    .S(net413),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _06982_ (.A0(net712),
    .A1(net1958),
    .S(net413),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _06983_ (.A0(net710),
    .A1(net1824),
    .S(net413),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _06984_ (.A0(net708),
    .A1(net2584),
    .S(net413),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _06985_ (.A0(net706),
    .A1(net2252),
    .S(net413),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _06986_ (.A0(net705),
    .A1(net1640),
    .S(net413),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _06987_ (.A0(net703),
    .A1(net2830),
    .S(net413),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _06988_ (.A0(net700),
    .A1(net2102),
    .S(net413),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _06989_ (.A0(net698),
    .A1(net2432),
    .S(net413),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _06990_ (.A0(net697),
    .A1(net2966),
    .S(net413),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _06991_ (.A0(net694),
    .A1(net2200),
    .S(net413),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _06992_ (.A0(net693),
    .A1(net2210),
    .S(net413),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _06993_ (.A0(net690),
    .A1(net2224),
    .S(net413),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _06994_ (.A0(net688),
    .A1(net2446),
    .S(net413),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _06995_ (.A0(net686),
    .A1(net1930),
    .S(net414),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _06996_ (.A0(net684),
    .A1(net2156),
    .S(net414),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _06997_ (.A0(net682),
    .A1(net2696),
    .S(net414),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _06998_ (.A0(net681),
    .A1(net2132),
    .S(net414),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _06999_ (.A0(net677),
    .A1(net2926),
    .S(net414),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _07000_ (.A0(net676),
    .A1(net2390),
    .S(net414),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _07001_ (.A0(net674),
    .A1(net2656),
    .S(net414),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _07002_ (.A0(net671),
    .A1(net1762),
    .S(net414),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _07003_ (.A0(net669),
    .A1(net2376),
    .S(net414),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _07004_ (.A0(net666),
    .A1(net1656),
    .S(net414),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _07005_ (.A0(net665),
    .A1(net3088),
    .S(net414),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _07006_ (.A0(net662),
    .A1(net3130),
    .S(net414),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _07007_ (.A0(net661),
    .A1(net2848),
    .S(net414),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _07008_ (.A0(net658),
    .A1(net1896),
    .S(net414),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _07009_ (.A0(net657),
    .A1(net1914),
    .S(net414),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _07010_ (.A0(net654),
    .A1(net2304),
    .S(net414),
    .X(_00041_));
 sky130_fd_sc_hd__or3_4 _07011_ (.A(\ctrl.c2d_rf_waddr_W[0] ),
    .B(_01777_),
    .C(_01818_),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_4 _07012_ (.A(_01808_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__mux2_1 _07013_ (.A0(net2864),
    .A1(net718),
    .S(net455),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _07014_ (.A0(net1650),
    .A1(net717),
    .S(net455),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _07015_ (.A0(net1754),
    .A1(net715),
    .S(net455),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _07016_ (.A0(net2320),
    .A1(net713),
    .S(net455),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _07017_ (.A0(net1704),
    .A1(net710),
    .S(net455),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _07018_ (.A0(net1920),
    .A1(net708),
    .S(net455),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _07019_ (.A0(net1924),
    .A1(net706),
    .S(net455),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _07020_ (.A0(net3040),
    .A1(net705),
    .S(net455),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _07021_ (.A0(net1800),
    .A1(net703),
    .S(net455),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _07022_ (.A0(net2596),
    .A1(net700),
    .S(net455),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _07023_ (.A0(net1984),
    .A1(net698),
    .S(net455),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _07024_ (.A0(net1582),
    .A1(net697),
    .S(net455),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _07025_ (.A0(net2774),
    .A1(net694),
    .S(net455),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _07026_ (.A0(net2916),
    .A1(net693),
    .S(net455),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _07027_ (.A0(net2464),
    .A1(net690),
    .S(net455),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _07028_ (.A0(net2664),
    .A1(net688),
    .S(net455),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _07029_ (.A0(net2196),
    .A1(net686),
    .S(net456),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _07030_ (.A0(net2894),
    .A1(net684),
    .S(net456),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _07031_ (.A0(net1558),
    .A1(net682),
    .S(net456),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _07032_ (.A0(net1460),
    .A1(net681),
    .S(net456),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _07033_ (.A0(net1554),
    .A1(net677),
    .S(net456),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _07034_ (.A0(net1292),
    .A1(net675),
    .S(net456),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(net2172),
    .A1(net673),
    .S(net456),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _07036_ (.A0(net1580),
    .A1(net671),
    .S(net456),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _07037_ (.A0(net2234),
    .A1(net668),
    .S(net456),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _07038_ (.A0(net1634),
    .A1(net666),
    .S(net456),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _07039_ (.A0(net2552),
    .A1(net665),
    .S(net456),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _07040_ (.A0(net2582),
    .A1(net662),
    .S(net456),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _07041_ (.A0(net2034),
    .A1(net661),
    .S(net456),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _07042_ (.A0(net1840),
    .A1(net658),
    .S(net456),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _07043_ (.A0(net2940),
    .A1(net657),
    .S(net456),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _07044_ (.A0(net1766),
    .A1(net654),
    .S(net456),
    .X(_00073_));
 sky130_fd_sc_hd__or4_4 _07045_ (.A(\ctrl.c2d_rf_waddr_W[0] ),
    .B(\ctrl.c2d_rf_waddr_W[1] ),
    .C(_01808_),
    .D(_01818_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _07046_ (.A0(net718),
    .A1(net2998),
    .S(net463),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(net717),
    .A1(net2548),
    .S(net463),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _07048_ (.A0(net714),
    .A1(net2944),
    .S(net463),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _07049_ (.A0(net712),
    .A1(net3070),
    .S(net463),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _07050_ (.A0(net710),
    .A1(net2646),
    .S(net463),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _07051_ (.A0(net708),
    .A1(net2384),
    .S(net463),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _07052_ (.A0(net706),
    .A1(net2892),
    .S(net463),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _07053_ (.A0(net705),
    .A1(net2784),
    .S(net463),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _07054_ (.A0(net703),
    .A1(net2002),
    .S(net463),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _07055_ (.A0(net700),
    .A1(net2734),
    .S(net463),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _07056_ (.A0(net698),
    .A1(net2316),
    .S(net463),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _07057_ (.A0(net697),
    .A1(net2718),
    .S(net463),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _07058_ (.A0(net694),
    .A1(net3074),
    .S(net463),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _07059_ (.A0(net693),
    .A1(net2094),
    .S(net463),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _07060_ (.A0(net690),
    .A1(net2754),
    .S(net463),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _07061_ (.A0(net688),
    .A1(net2640),
    .S(net463),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _07062_ (.A0(net686),
    .A1(net2684),
    .S(net464),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _07063_ (.A0(net684),
    .A1(net2618),
    .S(net464),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _07064_ (.A0(net682),
    .A1(net2986),
    .S(net464),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _07065_ (.A0(net681),
    .A1(net2182),
    .S(net464),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _07066_ (.A0(net677),
    .A1(net2282),
    .S(net464),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _07067_ (.A0(net675),
    .A1(net2276),
    .S(net464),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _07068_ (.A0(net673),
    .A1(net1940),
    .S(net464),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _07069_ (.A0(net671),
    .A1(net3048),
    .S(net464),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _07070_ (.A0(net669),
    .A1(net2788),
    .S(net464),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _07071_ (.A0(net666),
    .A1(net3150),
    .S(net464),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _07072_ (.A0(net665),
    .A1(net3192),
    .S(net464),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _07073_ (.A0(net662),
    .A1(net2232),
    .S(net464),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _07074_ (.A0(net661),
    .A1(net2244),
    .S(net464),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _07075_ (.A0(net658),
    .A1(net2808),
    .S(net464),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _07076_ (.A0(net657),
    .A1(net2764),
    .S(net464),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _07077_ (.A0(net654),
    .A1(net2712),
    .S(net464),
    .X(_00105_));
 sky130_fd_sc_hd__and3_2 _07078_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(\ctrl.c2d_rf_waddr_W[3] ),
    .C(\ctrl.c2d_rf_waddr_W[4] ),
    .X(_01826_));
 sky130_fd_sc_hd__or3_2 _07079_ (.A(_01778_),
    .B(_01779_),
    .C(_01780_),
    .X(_01827_));
 sky130_fd_sc_hd__nand2_4 _07080_ (.A(_01820_),
    .B(_01826_),
    .Y(_01828_));
 sky130_fd_sc_hd__mux2_1 _07081_ (.A0(net719),
    .A1(net2744),
    .S(net411),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _07082_ (.A0(net716),
    .A1(net2486),
    .S(net411),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _07083_ (.A0(net715),
    .A1(net3010),
    .S(net411),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _07084_ (.A0(net713),
    .A1(net3082),
    .S(net411),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _07085_ (.A0(net711),
    .A1(net2458),
    .S(net411),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _07086_ (.A0(net709),
    .A1(net3104),
    .S(net411),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _07087_ (.A0(net707),
    .A1(net3042),
    .S(net411),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _07088_ (.A0(net704),
    .A1(net2952),
    .S(net411),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _07089_ (.A0(net702),
    .A1(net3182),
    .S(net411),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _07090_ (.A0(net701),
    .A1(net2958),
    .S(net411),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _07091_ (.A0(net699),
    .A1(net2624),
    .S(net411),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _07092_ (.A0(net696),
    .A1(net3168),
    .S(net411),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _07093_ (.A0(net695),
    .A1(net2990),
    .S(net411),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _07094_ (.A0(net692),
    .A1(net2954),
    .S(net411),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _07095_ (.A0(net691),
    .A1(net2976),
    .S(net411),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _07096_ (.A0(net689),
    .A1(net2576),
    .S(net411),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _07097_ (.A0(net687),
    .A1(net2444),
    .S(net412),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _07098_ (.A0(net685),
    .A1(net2688),
    .S(net412),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _07099_ (.A0(net683),
    .A1(net2562),
    .S(net412),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _07100_ (.A0(net680),
    .A1(net2836),
    .S(net412),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _07101_ (.A0(net678),
    .A1(net2770),
    .S(net412),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _07102_ (.A0(net675),
    .A1(net2594),
    .S(net412),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _07103_ (.A0(net674),
    .A1(net3080),
    .S(net412),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _07104_ (.A0(net672),
    .A1(net2638),
    .S(net412),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _07105_ (.A0(net668),
    .A1(net3012),
    .S(net412),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _07106_ (.A0(net667),
    .A1(net3174),
    .S(net412),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _07107_ (.A0(net664),
    .A1(net3106),
    .S(net412),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _07108_ (.A0(net662),
    .A1(net3144),
    .S(net412),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _07109_ (.A0(net660),
    .A1(net3030),
    .S(net412),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _07110_ (.A0(\dpath.RF.wdata[29] ),
    .A1(net2702),
    .S(net412),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _07111_ (.A0(net656),
    .A1(net3076),
    .S(net412),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _07112_ (.A0(net654),
    .A1(net2898),
    .S(net412),
    .X(_00137_));
 sky130_fd_sc_hd__nor2_2 _07113_ (.A(\ctrl.c2d_rf_waddr_W[1] ),
    .B(_01819_),
    .Y(_01829_));
 sky130_fd_sc_hd__or2_4 _07114_ (.A(\ctrl.c2d_rf_waddr_W[1] ),
    .B(_01819_),
    .X(_01830_));
 sky130_fd_sc_hd__nand2_4 _07115_ (.A(_01826_),
    .B(_01829_),
    .Y(_01831_));
 sky130_fd_sc_hd__mux2_1 _07116_ (.A0(net719),
    .A1(net3180),
    .S(net409),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _07117_ (.A0(net716),
    .A1(net2612),
    .S(net409),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _07118_ (.A0(net715),
    .A1(net1870),
    .S(net409),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _07119_ (.A0(net713),
    .A1(net2900),
    .S(net409),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _07120_ (.A0(net711),
    .A1(net2628),
    .S(net409),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _07121_ (.A0(net709),
    .A1(net2700),
    .S(net409),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _07122_ (.A0(net707),
    .A1(net2606),
    .S(net409),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _07123_ (.A0(net704),
    .A1(net3028),
    .S(net409),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _07124_ (.A0(net702),
    .A1(net2920),
    .S(net409),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _07125_ (.A0(net701),
    .A1(net2874),
    .S(net409),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _07126_ (.A0(net699),
    .A1(net2970),
    .S(net409),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _07127_ (.A0(net696),
    .A1(net3172),
    .S(net409),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _07128_ (.A0(net695),
    .A1(net3102),
    .S(net409),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _07129_ (.A0(net692),
    .A1(net3140),
    .S(net409),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _07130_ (.A0(net691),
    .A1(net3126),
    .S(net409),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _07131_ (.A0(net689),
    .A1(net2914),
    .S(net409),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _07132_ (.A0(net687),
    .A1(net3078),
    .S(net410),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _07133_ (.A0(net685),
    .A1(net3020),
    .S(net410),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _07134_ (.A0(net683),
    .A1(net3124),
    .S(net410),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _07135_ (.A0(net680),
    .A1(net2978),
    .S(net410),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _07136_ (.A0(net678),
    .A1(net2710),
    .S(net410),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _07137_ (.A0(net675),
    .A1(net2984),
    .S(net410),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _07138_ (.A0(net674),
    .A1(net2194),
    .S(net410),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _07139_ (.A0(net672),
    .A1(net2860),
    .S(net410),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _07140_ (.A0(net668),
    .A1(net2572),
    .S(net410),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _07141_ (.A0(net667),
    .A1(net2616),
    .S(net410),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _07142_ (.A0(net664),
    .A1(net2466),
    .S(net410),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _07143_ (.A0(net662),
    .A1(net3128),
    .S(net410),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _07144_ (.A0(net660),
    .A1(net2852),
    .S(net410),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _07145_ (.A0(net658),
    .A1(net2636),
    .S(net410),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _07146_ (.A0(net656),
    .A1(net2374),
    .S(net410),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _07147_ (.A0(net654),
    .A1(net2238),
    .S(net410),
    .X(_00169_));
 sky130_fd_sc_hd__or3_4 _07148_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(\ctrl.c2d_rf_waddr_W[3] ),
    .C(\ctrl.c2d_rf_waddr_W[4] ),
    .X(_01832_));
 sky130_fd_sc_hd__or2_4 _07149_ (.A(_01821_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _07150_ (.A0(net718),
    .A1(net3152),
    .S(net407),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _07151_ (.A0(net717),
    .A1(net2838),
    .S(net407),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _07152_ (.A0(net714),
    .A1(net2442),
    .S(net407),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _07153_ (.A0(net712),
    .A1(net2420),
    .S(net407),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _07154_ (.A0(net710),
    .A1(net2814),
    .S(net407),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _07155_ (.A0(net708),
    .A1(net3118),
    .S(net407),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _07156_ (.A0(net706),
    .A1(net3186),
    .S(net407),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _07157_ (.A0(net705),
    .A1(net2354),
    .S(net407),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _07158_ (.A0(net702),
    .A1(net2644),
    .S(net407),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _07159_ (.A0(net700),
    .A1(net2796),
    .S(net407),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _07160_ (.A0(net698),
    .A1(net2418),
    .S(net407),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _07161_ (.A0(net697),
    .A1(net2794),
    .S(net407),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _07162_ (.A0(net695),
    .A1(net2256),
    .S(net407),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _07163_ (.A0(net693),
    .A1(net2508),
    .S(net407),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _07164_ (.A0(net690),
    .A1(net1968),
    .S(net407),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _07165_ (.A0(net688),
    .A1(net2214),
    .S(net407),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _07166_ (.A0(net686),
    .A1(net2974),
    .S(net408),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _07167_ (.A0(net684),
    .A1(net2522),
    .S(net408),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _07168_ (.A0(net682),
    .A1(net2742),
    .S(net408),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _07169_ (.A0(net681),
    .A1(net2896),
    .S(net408),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _07170_ (.A0(net677),
    .A1(net3120),
    .S(net408),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _07171_ (.A0(net676),
    .A1(net2670),
    .S(net408),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _07172_ (.A0(net673),
    .A1(net2558),
    .S(net408),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _07173_ (.A0(net671),
    .A1(net2750),
    .S(net408),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _07174_ (.A0(net669),
    .A1(net2534),
    .S(net408),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _07175_ (.A0(net666),
    .A1(net2768),
    .S(net408),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _07176_ (.A0(net665),
    .A1(net2674),
    .S(net408),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _07177_ (.A0(net662),
    .A1(net2072),
    .S(net408),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _07178_ (.A0(net661),
    .A1(net2298),
    .S(net408),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _07179_ (.A0(net659),
    .A1(net2826),
    .S(net408),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _07180_ (.A0(net657),
    .A1(net2402),
    .S(net408),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _07181_ (.A0(net654),
    .A1(net2510),
    .S(net408),
    .X(_00201_));
 sky130_fd_sc_hd__nor2_4 _07182_ (.A(_01808_),
    .B(_01830_),
    .Y(_01834_));
 sky130_fd_sc_hd__mux2_1 _07183_ (.A0(net2932),
    .A1(net718),
    .S(net405),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _07184_ (.A0(net2542),
    .A1(net717),
    .S(net405),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _07185_ (.A0(net1996),
    .A1(net714),
    .S(net405),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _07186_ (.A0(net1576),
    .A1(net712),
    .S(net405),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _07187_ (.A0(net2048),
    .A1(net710),
    .S(net405),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _07188_ (.A0(net1282),
    .A1(net708),
    .S(net405),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _07189_ (.A0(net2782),
    .A1(net706),
    .S(net405),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _07190_ (.A0(net1612),
    .A1(net705),
    .S(net405),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _07191_ (.A0(net1316),
    .A1(net703),
    .S(net405),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _07192_ (.A0(net2600),
    .A1(net700),
    .S(net405),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _07193_ (.A0(net2720),
    .A1(net698),
    .S(net405),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _07194_ (.A0(net1786),
    .A1(net697),
    .S(net405),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _07195_ (.A0(net1198),
    .A1(net694),
    .S(net405),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _07196_ (.A0(net2866),
    .A1(net693),
    .S(net405),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _07197_ (.A0(net2748),
    .A1(net690),
    .S(net405),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _07198_ (.A0(net1608),
    .A1(net688),
    .S(net405),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _07199_ (.A0(net2338),
    .A1(net686),
    .S(net406),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _07200_ (.A0(net1186),
    .A1(net684),
    .S(net406),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _07201_ (.A0(net1950),
    .A1(net682),
    .S(net406),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _07202_ (.A0(net2330),
    .A1(net681),
    .S(net406),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _07203_ (.A0(net1512),
    .A1(net677),
    .S(net406),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _07204_ (.A0(net1516),
    .A1(net676),
    .S(net406),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _07205_ (.A0(net1570),
    .A1(net673),
    .S(net406),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _07206_ (.A0(net1734),
    .A1(net671),
    .S(net406),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _07207_ (.A0(net2030),
    .A1(net668),
    .S(net406),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _07208_ (.A0(net2398),
    .A1(net667),
    .S(net406),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _07209_ (.A0(net3166),
    .A1(net665),
    .S(net406),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _07210_ (.A0(net1670),
    .A1(net663),
    .S(net406),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _07211_ (.A0(net1188),
    .A1(net661),
    .S(net406),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _07212_ (.A0(net2346),
    .A1(net658),
    .S(net406),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _07213_ (.A0(net1296),
    .A1(net657),
    .S(net406),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _07214_ (.A0(net2042),
    .A1(net655),
    .S(net406),
    .X(_00233_));
 sky130_fd_sc_hd__and4b_1 _07215_ (.A_N(\ctrl.d2c_inst[4] ),
    .B(\ctrl.d2c_inst[1] ),
    .C(\ctrl.d2c_inst[0] ),
    .D(\ctrl.d2c_inst[5] ),
    .X(_01835_));
 sky130_fd_sc_hd__and4_4 _07216_ (.A(net3345),
    .B(net3176),
    .C(net3211),
    .D(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__or4bb_2 _07217_ (.A(net1150),
    .B(\ctrl.inst_X[2] ),
    .C_N(\ctrl.inst_X[1] ),
    .D_N(\ctrl.inst_X[0] ),
    .X(_01837_));
 sky130_fd_sc_hd__and3b_1 _07218_ (.A_N(\ctrl.inst_X[4] ),
    .B(\ctrl.inst_X[5] ),
    .C(\ctrl.inst_X[6] ),
    .X(_01838_));
 sky130_fd_sc_hd__nor2_1 _07219_ (.A(\ctrl.inst_X[14] ),
    .B(\ctrl.inst_X[13] ),
    .Y(_01839_));
 sky130_fd_sc_hd__or4bb_2 _07220_ (.A(_01763_),
    .B(_01837_),
    .C_N(_01838_),
    .D_N(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__and2_1 _07222_ (.A(net651),
    .B(net786),
    .X(_01842_));
 sky130_fd_sc_hd__nor2_1 _07223_ (.A(net651),
    .B(net786),
    .Y(_01843_));
 sky130_fd_sc_hd__nor2_1 _07224_ (.A(_01842_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__and2_2 _07225_ (.A(net628),
    .B(net768),
    .X(_01845_));
 sky130_fd_sc_hd__nor2_1 _07226_ (.A(\dpath.alu.adder.in0[5] ),
    .B(net768),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _07227_ (.A(_01845_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(net601),
    .B(net742),
    .Y(_01848_));
 sky130_fd_sc_hd__or2_1 _07229_ (.A(net601),
    .B(net742),
    .X(_01849_));
 sky130_fd_sc_hd__and2_1 _07230_ (.A(_01848_),
    .B(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__and2_1 _07231_ (.A(\dpath.alu.adder.in0[4] ),
    .B(net772),
    .X(_01851_));
 sky130_fd_sc_hd__nor2_1 _07232_ (.A(\dpath.alu.adder.in0[4] ),
    .B(net772),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _07233_ (.A(_01851_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_2 _07234_ (.A(net643),
    .B(net780),
    .Y(_01854_));
 sky130_fd_sc_hd__inv_2 _07235_ (.A(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _07236_ (.A(net643),
    .B(net780),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _07237_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__or2_1 _07238_ (.A(\dpath.alu.adder.in0[29] ),
    .B(\dpath.alu.adder.in1[29] ),
    .X(_01858_));
 sky130_fd_sc_hd__nand2_1 _07239_ (.A(\dpath.alu.adder.in0[29] ),
    .B(\dpath.alu.adder.in1[29] ),
    .Y(_01859_));
 sky130_fd_sc_hd__and2_1 _07240_ (.A(_01858_),
    .B(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__nor2_1 _07241_ (.A(net590),
    .B(net731),
    .Y(_01861_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(net590),
    .B(net730),
    .Y(_01862_));
 sky130_fd_sc_hd__and2b_1 _07243_ (.A_N(_01861_),
    .B(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__nand2_2 _07244_ (.A(net616),
    .B(net757),
    .Y(_01864_));
 sky130_fd_sc_hd__or2_1 _07245_ (.A(net616),
    .B(net757),
    .X(_01865_));
 sky130_fd_sc_hd__nand2_1 _07246_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand2_1 _07247_ (.A(net584),
    .B(net725),
    .Y(_01867_));
 sky130_fd_sc_hd__or2_1 _07248_ (.A(net583),
    .B(net725),
    .X(_01868_));
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__and2_1 _07250_ (.A(net613),
    .B(net754),
    .X(_01870_));
 sky130_fd_sc_hd__nor2_1 _07251_ (.A(net613),
    .B(net754),
    .Y(_01871_));
 sky130_fd_sc_hd__or2_1 _07252_ (.A(_01870_),
    .B(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__nor2_1 _07253_ (.A(\dpath.alu.adder.in0[27] ),
    .B(\dpath.alu.adder.in1[27] ),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _07254_ (.A(\dpath.alu.adder.in0[27] ),
    .B(\dpath.alu.adder.in1[27] ),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2b_2 _07255_ (.A_N(_01873_),
    .B(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(net604),
    .B(net746),
    .Y(_01876_));
 sky130_fd_sc_hd__or2_1 _07257_ (.A(net604),
    .B(net746),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_2 _07258_ (.A(_01876_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _07259_ (.A(net581),
    .B(net724),
    .Y(_01879_));
 sky130_fd_sc_hd__or2_1 _07260_ (.A(net581),
    .B(net724),
    .X(_01880_));
 sky130_fd_sc_hd__nand2_1 _07261_ (.A(_01879_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(\dpath.alu.adder.in0[30] ),
    .B(\dpath.alu.adder.in1[30] ),
    .Y(_01882_));
 sky130_fd_sc_hd__or2_1 _07263_ (.A(\dpath.alu.adder.in0[30] ),
    .B(\dpath.alu.adder.in1[30] ),
    .X(_01883_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(_01882_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_2 _07265_ (.A(net607),
    .B(net750),
    .Y(_01885_));
 sky130_fd_sc_hd__or2_1 _07266_ (.A(net607),
    .B(net750),
    .X(_01886_));
 sky130_fd_sc_hd__and2_1 _07267_ (.A(_01885_),
    .B(_01886_),
    .X(_01887_));
 sky130_fd_sc_hd__inv_2 _07268_ (.A(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__or2_1 _07269_ (.A(net592),
    .B(net732),
    .X(_01889_));
 sky130_fd_sc_hd__nand2_1 _07270_ (.A(net592),
    .B(net732),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _07271_ (.A(_01889_),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__or2_1 _07272_ (.A(\dpath.alu.adder.in0[25] ),
    .B(\dpath.alu.adder.in1[25] ),
    .X(_01892_));
 sky130_fd_sc_hd__nand2_1 _07273_ (.A(\dpath.alu.adder.in0[25] ),
    .B(\dpath.alu.adder.in1[25] ),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_2 _07274_ (.A(_01892_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand2_2 _07275_ (.A(net598),
    .B(net736),
    .Y(_01895_));
 sky130_fd_sc_hd__or2_1 _07276_ (.A(net598),
    .B(net736),
    .X(_01896_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(_01895_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__or2_1 _07278_ (.A(\dpath.alu.adder.in0[24] ),
    .B(\dpath.alu.adder.in1[24] ),
    .X(_01898_));
 sky130_fd_sc_hd__nand2_1 _07279_ (.A(\dpath.alu.adder.in0[24] ),
    .B(\dpath.alu.adder.in1[24] ),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(_01898_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__or2_1 _07281_ (.A(net638),
    .B(net776),
    .X(_01901_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(net638),
    .B(net776),
    .Y(_01902_));
 sky130_fd_sc_hd__nand2_1 _07283_ (.A(_01901_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__and2_1 _07284_ (.A(net647),
    .B(net783),
    .X(_01904_));
 sky130_fd_sc_hd__xor2_2 _07285_ (.A(net647),
    .B(net783),
    .X(_01905_));
 sky130_fd_sc_hd__xor2_2 _07286_ (.A(\dpath.alu.adder.in0[31] ),
    .B(\dpath.alu.adder.in1[31] ),
    .X(_01906_));
 sky130_fd_sc_hd__inv_2 _07287_ (.A(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _07288_ (.A(net596),
    .B(net734),
    .Y(_01908_));
 sky130_fd_sc_hd__or2_1 _07289_ (.A(net595),
    .B(net734),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _07290_ (.A(_01908_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand2_1 _07291_ (.A(net585),
    .B(net727),
    .Y(_01911_));
 sky130_fd_sc_hd__or2_1 _07292_ (.A(net585),
    .B(net727),
    .X(_01912_));
 sky130_fd_sc_hd__nand2_1 _07293_ (.A(_01911_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__or2_1 _07294_ (.A(\dpath.alu.adder.in0[26] ),
    .B(\dpath.alu.adder.in1[26] ),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_1 _07295_ (.A(\dpath.alu.adder.in0[26] ),
    .B(net3635),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _07296_ (.A(_01914_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _07297_ (.A(net579),
    .B(\dpath.alu.adder.in1[23] ),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(net579),
    .B(net721),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2b_1 _07299_ (.A_N(_01917_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__or2_1 _07300_ (.A(\dpath.alu.adder.in0[22] ),
    .B(net722),
    .X(_01920_));
 sky130_fd_sc_hd__nand2_2 _07301_ (.A(\dpath.alu.adder.in0[22] ),
    .B(\dpath.alu.adder.in1[22] ),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_2 _07302_ (.A(_01920_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__and2_1 _07303_ (.A(net611),
    .B(net751),
    .X(_01923_));
 sky130_fd_sc_hd__nor2_1 _07304_ (.A(net611),
    .B(net751),
    .Y(_01924_));
 sky130_fd_sc_hd__nor2_1 _07305_ (.A(_01923_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _07306_ (.A(net624),
    .B(net764),
    .Y(_01926_));
 sky130_fd_sc_hd__or2_1 _07307_ (.A(net624),
    .B(net764),
    .X(_01927_));
 sky130_fd_sc_hd__nand2_1 _07308_ (.A(_01926_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__inv_2 _07309_ (.A(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_1 _07310_ (.A(net587),
    .B(net729),
    .Y(_01930_));
 sky130_fd_sc_hd__or2_1 _07311_ (.A(net587),
    .B(net729),
    .X(_01931_));
 sky130_fd_sc_hd__nand2_1 _07312_ (.A(_01930_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__and2_1 _07313_ (.A(net620),
    .B(net760),
    .X(_01933_));
 sky130_fd_sc_hd__or2_1 _07314_ (.A(net620),
    .B(net760),
    .X(_01934_));
 sky130_fd_sc_hd__nand2b_1 _07315_ (.A_N(_01933_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__or2_1 _07316_ (.A(\dpath.alu.adder.in0[28] ),
    .B(\dpath.alu.adder.in1[28] ),
    .X(_01936_));
 sky130_fd_sc_hd__nand2_1 _07317_ (.A(\dpath.alu.adder.in0[28] ),
    .B(\dpath.alu.adder.in1[28] ),
    .Y(_01937_));
 sky130_fd_sc_hd__and2_1 _07318_ (.A(_01936_),
    .B(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__and4_1 _07319_ (.A(_01866_),
    .B(_01872_),
    .C(_01875_),
    .D(_01922_),
    .X(_01939_));
 sky130_fd_sc_hd__and4_1 _07320_ (.A(_01869_),
    .B(_01878_),
    .C(_01881_),
    .D(_01919_),
    .X(_01940_));
 sky130_fd_sc_hd__nand3_1 _07321_ (.A(_01841_),
    .B(_01939_),
    .C(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand3_1 _07322_ (.A(_01900_),
    .B(_01910_),
    .C(_01916_),
    .Y(_01942_));
 sky130_fd_sc_hd__or4_1 _07323_ (.A(_01844_),
    .B(_01850_),
    .C(_01853_),
    .D(_01857_),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_1 _07324_ (.A(_01928_),
    .B(_01935_),
    .Y(_01944_));
 sky130_fd_sc_hd__or4b_1 _07325_ (.A(_01860_),
    .B(_01863_),
    .C(_01925_),
    .D_N(_01932_),
    .X(_01945_));
 sky130_fd_sc_hd__or4_1 _07326_ (.A(_01906_),
    .B(_01938_),
    .C(_01944_),
    .D(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__nand3_1 _07327_ (.A(_01894_),
    .B(_01897_),
    .C(_01903_),
    .Y(_01947_));
 sky130_fd_sc_hd__and4_1 _07328_ (.A(_01884_),
    .B(_01888_),
    .C(_01891_),
    .D(_01913_),
    .X(_01948_));
 sky130_fd_sc_hd__or4b_1 _07329_ (.A(_01905_),
    .B(_01946_),
    .C(_01947_),
    .D_N(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__or4_1 _07330_ (.A(_01847_),
    .B(_01942_),
    .C(_01943_),
    .D(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__o2bb2a_1 _07331_ (.A1_N(_01840_),
    .A2_N(_01844_),
    .B1(_01941_),
    .B2(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__and3_4 _07332_ (.A(net3327),
    .B(_01841_),
    .C(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__and4bb_1 _07333_ (.A_N(\ctrl.d2c_inst[12] ),
    .B_N(\ctrl.d2c_inst[3] ),
    .C(\ctrl.d2c_inst[2] ),
    .D(\ctrl.d2c_inst[6] ),
    .X(_01953_));
 sky130_fd_sc_hd__and4bb_1 _07334_ (.A_N(net3715),
    .B_N(net3282),
    .C(_01835_),
    .D(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__nand2_1 _07335_ (.A(net3465),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2b_1 _07336_ (.A_N(net404),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__a21oi_1 _07337_ (.A1(net3465),
    .A2(_01836_),
    .B1(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__a21o_4 _07338_ (.A1(net3465),
    .A2(_01836_),
    .B1(_01956_),
    .X(_01958_));
 sky130_fd_sc_hd__nor3_1 _07339_ (.A(\ctrl.inst_X[6] ),
    .B(\ctrl.inst_X[12] ),
    .C(_01837_),
    .Y(_01959_));
 sky130_fd_sc_hd__inv_2 _07340_ (.A(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__or4b_4 _07341_ (.A(net3207),
    .B(_01960_),
    .C(net2972),
    .D_N(net2868),
    .X(_01961_));
 sky130_fd_sc_hd__or2_1 _07342_ (.A(\ctrl.inst_X[5] ),
    .B(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__or4_1 _07343_ (.A(\ctrl.inst_X[7] ),
    .B(\ctrl.inst_X[8] ),
    .C(\ctrl.inst_X[10] ),
    .D(\ctrl.inst_X[11] ),
    .X(_01963_));
 sky130_fd_sc_hd__o21ba_1 _07344_ (.A1(net3245),
    .A2(_01963_),
    .B1_N(_01962_),
    .X(_01964_));
 sky130_fd_sc_hd__or4bb_2 _07345_ (.A(net3531),
    .B(net3276),
    .C_N(\ctrl.d2c_inst[1] ),
    .D_N(\ctrl.d2c_inst[0] ),
    .X(_01965_));
 sky130_fd_sc_hd__or2_1 _07346_ (.A(net3470),
    .B(\ctrl.d2c_inst[6] ),
    .X(_01966_));
 sky130_fd_sc_hd__or2_1 _07347_ (.A(_01965_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__or4_1 _07348_ (.A(\ctrl.d2c_inst[29] ),
    .B(\ctrl.d2c_inst[28] ),
    .C(\ctrl.d2c_inst[27] ),
    .D(\ctrl.d2c_inst[26] ),
    .X(_01968_));
 sky130_fd_sc_hd__nand2_1 _07349_ (.A(net3499),
    .B(\ctrl.d2c_inst[4] ),
    .Y(_01969_));
 sky130_fd_sc_hd__or4_1 _07350_ (.A(net577),
    .B(\ctrl.d2c_inst[30] ),
    .C(\ctrl.d2c_inst[14] ),
    .D(\ctrl.d2c_inst[13] ),
    .X(_01970_));
 sky130_fd_sc_hd__nor4_1 _07351_ (.A(_01967_),
    .B(_01968_),
    .C(_01969_),
    .D(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__and4bb_1 _07352_ (.A_N(\ctrl.d2c_inst[14] ),
    .B_N(\ctrl.d2c_inst[13] ),
    .C(\ctrl.d2c_inst[12] ),
    .D(\ctrl.d2c_inst[6] ),
    .X(_01972_));
 sky130_fd_sc_hd__and4bb_2 _07353_ (.A_N(net3550),
    .B_N(_01965_),
    .C(_01972_),
    .D(net3499),
    .X(_01973_));
 sky130_fd_sc_hd__or4b_2 _07354_ (.A(_01759_),
    .B(net3429),
    .C(_01965_),
    .D_N(_01972_),
    .X(_01974_));
 sky130_fd_sc_hd__nor2_4 _07355_ (.A(net481),
    .B(_01973_),
    .Y(_01975_));
 sky130_fd_sc_hd__or3b_1 _07356_ (.A(\ctrl.d2c_inst[14] ),
    .B(\ctrl.d2c_inst[4] ),
    .C_N(\ctrl.d2c_inst[13] ),
    .X(_01976_));
 sky130_fd_sc_hd__or4b_1 _07357_ (.A(\ctrl.d2c_inst[14] ),
    .B(\ctrl.d2c_inst[13] ),
    .C(\ctrl.d2c_inst[5] ),
    .D_N(\ctrl.d2c_inst[4] ),
    .X(_01977_));
 sky130_fd_sc_hd__a21o_1 _07358_ (.A1(_01976_),
    .A2(_01977_),
    .B1(_01967_),
    .X(_01978_));
 sky130_fd_sc_hd__or4b_1 _07359_ (.A(_01954_),
    .B(_01971_),
    .C(_01973_),
    .D_N(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__nor3b_1 _07360_ (.A(_01965_),
    .B(_01969_),
    .C_N(_01972_),
    .Y(_01980_));
 sky130_fd_sc_hd__o21a_1 _07361_ (.A1(net475),
    .A2(_01980_),
    .B1(\ctrl.val_D ),
    .X(_01981_));
 sky130_fd_sc_hd__or4_4 _07362_ (.A(_01759_),
    .B(_01965_),
    .C(_01966_),
    .D(_01976_),
    .X(_01982_));
 sky130_fd_sc_hd__a21boi_2 _07363_ (.A1(net478),
    .A2(_01982_),
    .B1_N(\ctrl.val_D ),
    .Y(_01983_));
 sky130_fd_sc_hd__xor2_1 _07364_ (.A(\ctrl.d2c_inst[24] ),
    .B(\ctrl.inst_X[11] ),
    .X(_01984_));
 sky130_fd_sc_hd__or2_1 _07365_ (.A(\ctrl.d2c_inst[23] ),
    .B(\ctrl.inst_X[10] ),
    .X(_01985_));
 sky130_fd_sc_hd__nand2_1 _07366_ (.A(\ctrl.d2c_inst[23] ),
    .B(\ctrl.inst_X[10] ),
    .Y(_01986_));
 sky130_fd_sc_hd__or2_1 _07367_ (.A(\ctrl.d2c_inst[22] ),
    .B(\ctrl.inst_X[9] ),
    .X(_01987_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(\ctrl.d2c_inst[22] ),
    .B(\ctrl.inst_X[9] ),
    .Y(_01988_));
 sky130_fd_sc_hd__a22o_1 _07369_ (.A1(_01985_),
    .A2(_01986_),
    .B1(_01987_),
    .B2(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__or2_1 _07370_ (.A(\ctrl.d2c_inst[20] ),
    .B(\ctrl.inst_X[7] ),
    .X(_01990_));
 sky130_fd_sc_hd__nand2_1 _07371_ (.A(\ctrl.d2c_inst[20] ),
    .B(\ctrl.inst_X[7] ),
    .Y(_01991_));
 sky130_fd_sc_hd__or2_1 _07372_ (.A(\ctrl.d2c_inst[21] ),
    .B(\ctrl.inst_X[8] ),
    .X(_01992_));
 sky130_fd_sc_hd__nand2_1 _07373_ (.A(\ctrl.d2c_inst[21] ),
    .B(\ctrl.inst_X[8] ),
    .Y(_01993_));
 sky130_fd_sc_hd__a221o_1 _07374_ (.A1(_01990_),
    .A2(_01991_),
    .B1(_01992_),
    .B2(_01993_),
    .C1(_01989_),
    .X(_01994_));
 sky130_fd_sc_hd__and4bb_1 _07375_ (.A_N(_01984_),
    .B_N(_01994_),
    .C(\ctrl.val_DX.q ),
    .D(_01983_),
    .X(_01995_));
 sky130_fd_sc_hd__o22a_1 _07376_ (.A1(_01755_),
    .A2(\ctrl.inst_X[10] ),
    .B1(_01768_),
    .B2(\ctrl.d2c_inst[19] ),
    .X(_01996_));
 sky130_fd_sc_hd__o22a_1 _07377_ (.A1(_01758_),
    .A2(\ctrl.inst_X[7] ),
    .B1(_01766_),
    .B2(\ctrl.d2c_inst[17] ),
    .X(_01997_));
 sky130_fd_sc_hd__o221a_1 _07378_ (.A1(\ctrl.d2c_inst[16] ),
    .A2(_01765_),
    .B1(\ctrl.inst_X[9] ),
    .B2(_01756_),
    .C1(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__o221a_1 _07379_ (.A1(\ctrl.d2c_inst[15] ),
    .A2(_01764_),
    .B1(\ctrl.inst_X[11] ),
    .B2(_01754_),
    .C1(_01996_),
    .X(_01999_));
 sky130_fd_sc_hd__o221a_1 _07380_ (.A1(_01757_),
    .A2(\ctrl.inst_X[8] ),
    .B1(_01767_),
    .B2(\ctrl.d2c_inst[18] ),
    .C1(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__and4_2 _07381_ (.A(\ctrl.val_DX.q ),
    .B(_01981_),
    .C(_01998_),
    .D(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__o22a_1 _07382_ (.A1(_01750_),
    .A2(\ctrl.inst_X[10] ),
    .B1(_01768_),
    .B2(\ctrl.d2c_inst[24] ),
    .X(_02002_));
 sky130_fd_sc_hd__o22a_1 _07383_ (.A1(_01753_),
    .A2(\ctrl.inst_X[7] ),
    .B1(_01766_),
    .B2(\ctrl.d2c_inst[22] ),
    .X(_02003_));
 sky130_fd_sc_hd__o221a_1 _07384_ (.A1(\ctrl.d2c_inst[21] ),
    .A2(_01765_),
    .B1(\ctrl.inst_X[9] ),
    .B2(_01751_),
    .C1(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__o221a_1 _07385_ (.A1(\ctrl.d2c_inst[20] ),
    .A2(_01764_),
    .B1(\ctrl.inst_X[11] ),
    .B2(_01749_),
    .C1(_02002_),
    .X(_02005_));
 sky130_fd_sc_hd__o221a_1 _07386_ (.A1(_01752_),
    .A2(\ctrl.inst_X[8] ),
    .B1(_01767_),
    .B2(\ctrl.d2c_inst[23] ),
    .C1(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__and4_2 _07387_ (.A(\ctrl.val_DX.q ),
    .B(_01983_),
    .C(_02004_),
    .D(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__o21a_2 _07388_ (.A1(_02001_),
    .A2(_02007_),
    .B1(_01964_),
    .X(_02008_));
 sky130_fd_sc_hd__o21ai_4 _07389_ (.A1(_02001_),
    .A2(_02007_),
    .B1(_01964_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_2 _07390_ (.A(net362),
    .B(net452),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(_01958_),
    .B(net446),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _07392_ (.A(net880),
    .B(_02010_),
    .Y(_00234_));
 sky130_fd_sc_hd__and2_1 _07393_ (.A(net3198),
    .B(net857),
    .X(_00235_));
 sky130_fd_sc_hd__and2_1 _07394_ (.A(net1176),
    .B(net854),
    .X(_00236_));
 sky130_fd_sc_hd__and2_1 _07395_ (.A(net1208),
    .B(net854),
    .X(_00237_));
 sky130_fd_sc_hd__and2_1 _07396_ (.A(net1166),
    .B(net854),
    .X(_00238_));
 sky130_fd_sc_hd__and2_1 _07397_ (.A(net1150),
    .B(net854),
    .X(_00239_));
 sky130_fd_sc_hd__and2_1 _07398_ (.A(net3207),
    .B(net855),
    .X(_00240_));
 sky130_fd_sc_hd__and2_1 _07399_ (.A(net3209),
    .B(net856),
    .X(_00241_));
 sky130_fd_sc_hd__and2_1 _07400_ (.A(net1468),
    .B(net855),
    .X(_00242_));
 sky130_fd_sc_hd__nor2_1 _07401_ (.A(_01764_),
    .B(net890),
    .Y(_00243_));
 sky130_fd_sc_hd__nor2_1 _07402_ (.A(_01765_),
    .B(net890),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_1 _07403_ (.A(_01766_),
    .B(net890),
    .Y(_00245_));
 sky130_fd_sc_hd__nor2_1 _07404_ (.A(_01767_),
    .B(net890),
    .Y(_00246_));
 sky130_fd_sc_hd__nor2_1 _07405_ (.A(_01768_),
    .B(net890),
    .Y(_00247_));
 sky130_fd_sc_hd__nor2_1 _07406_ (.A(net1157),
    .B(net893),
    .Y(_00248_));
 sky130_fd_sc_hd__and2_1 _07407_ (.A(net2868),
    .B(net855),
    .X(_00249_));
 sky130_fd_sc_hd__and2_1 _07408_ (.A(net2972),
    .B(net855),
    .X(_00250_));
 sky130_fd_sc_hd__and2_1 _07409_ (.A(net876),
    .B(net3436),
    .X(_00251_));
 sky130_fd_sc_hd__and2_1 _07410_ (.A(net876),
    .B(net3307),
    .X(_00252_));
 sky130_fd_sc_hd__and2_1 _07411_ (.A(net876),
    .B(net3424),
    .X(_00253_));
 sky130_fd_sc_hd__and2_1 _07412_ (.A(net876),
    .B(net3312),
    .X(_00254_));
 sky130_fd_sc_hd__and2_1 _07413_ (.A(net857),
    .B(net1000),
    .X(_00255_));
 sky130_fd_sc_hd__and2_1 _07414_ (.A(net1092),
    .B(net856),
    .X(_00256_));
 sky130_fd_sc_hd__and2_1 _07415_ (.A(net990),
    .B(net855),
    .X(_00257_));
 sky130_fd_sc_hd__and2_1 _07416_ (.A(net910),
    .B(net861),
    .X(_00258_));
 sky130_fd_sc_hd__and2_1 _07417_ (.A(net906),
    .B(net861),
    .X(_00259_));
 sky130_fd_sc_hd__and2_1 _07418_ (.A(net914),
    .B(net861),
    .X(_00260_));
 sky130_fd_sc_hd__and2_1 _07419_ (.A(net912),
    .B(net861),
    .X(_00261_));
 sky130_fd_sc_hd__and2_1 _07420_ (.A(net1090),
    .B(net856),
    .X(_00262_));
 sky130_fd_sc_hd__and4b_1 _07421_ (.A_N(net404),
    .B(net3465),
    .C(net854),
    .D(net446),
    .X(_00263_));
 sky130_fd_sc_hd__and2_1 _07422_ (.A(net2060),
    .B(net853),
    .X(_00264_));
 sky130_fd_sc_hd__and2_1 _07423_ (.A(net2406),
    .B(net853),
    .X(_00265_));
 sky130_fd_sc_hd__and2_1 _07424_ (.A(net3211),
    .B(net853),
    .X(_00266_));
 sky130_fd_sc_hd__and2_1 _07425_ (.A(net3176),
    .B(net853),
    .X(_00267_));
 sky130_fd_sc_hd__and2_1 _07426_ (.A(net3429),
    .B(net855),
    .X(_00268_));
 sky130_fd_sc_hd__nor2_1 _07427_ (.A(_01759_),
    .B(net893),
    .Y(_00269_));
 sky130_fd_sc_hd__and2_1 _07428_ (.A(net3345),
    .B(net853),
    .X(_00270_));
 sky130_fd_sc_hd__and2_1 _07429_ (.A(net3205),
    .B(net854),
    .X(_00271_));
 sky130_fd_sc_hd__and2_1 _07430_ (.A(net3235),
    .B(net855),
    .X(_00272_));
 sky130_fd_sc_hd__and2_1 _07431_ (.A(net3202),
    .B(net855),
    .X(_00273_));
 sky130_fd_sc_hd__and2_1 _07432_ (.A(net3237),
    .B(net854),
    .X(_00274_));
 sky130_fd_sc_hd__and2_1 _07433_ (.A(net3219),
    .B(net856),
    .X(_00275_));
 sky130_fd_sc_hd__and2_1 _07434_ (.A(net3264),
    .B(net855),
    .X(_00276_));
 sky130_fd_sc_hd__and2_1 _07435_ (.A(net3282),
    .B(net855),
    .X(_00277_));
 sky130_fd_sc_hd__and2_1 _07436_ (.A(net3342),
    .B(net855),
    .X(_00278_));
 sky130_fd_sc_hd__nor2_1 _07437_ (.A(_01753_),
    .B(net890),
    .Y(_00279_));
 sky130_fd_sc_hd__nor2_1 _07438_ (.A(_01752_),
    .B(net890),
    .Y(_00280_));
 sky130_fd_sc_hd__nor2_1 _07439_ (.A(_01751_),
    .B(net890),
    .Y(_00281_));
 sky130_fd_sc_hd__nor2_1 _07440_ (.A(_01750_),
    .B(net891),
    .Y(_00282_));
 sky130_fd_sc_hd__nor2_1 _07441_ (.A(_01749_),
    .B(net890),
    .Y(_00283_));
 sky130_fd_sc_hd__and2_1 _07442_ (.A(net3392),
    .B(net855),
    .X(_00284_));
 sky130_fd_sc_hd__and2_1 _07443_ (.A(net3452),
    .B(net860),
    .X(_00285_));
 sky130_fd_sc_hd__and2_1 _07444_ (.A(net3420),
    .B(net860),
    .X(_00286_));
 sky130_fd_sc_hd__and2_1 _07445_ (.A(net3421),
    .B(net860),
    .X(_00287_));
 sky130_fd_sc_hd__and2_1 _07446_ (.A(net3461),
    .B(net860),
    .X(_00288_));
 sky130_fd_sc_hd__and2_1 _07447_ (.A(net3435),
    .B(net860),
    .X(_00289_));
 sky130_fd_sc_hd__and2_1 _07448_ (.A(net3216),
    .B(net855),
    .X(_00290_));
 sky130_fd_sc_hd__and2_1 _07449_ (.A(net1022),
    .B(net854),
    .X(_00291_));
 sky130_fd_sc_hd__and2_1 _07450_ (.A(net972),
    .B(net854),
    .X(_00292_));
 sky130_fd_sc_hd__and2_1 _07451_ (.A(net3208),
    .B(net856),
    .X(_00293_));
 sky130_fd_sc_hd__and2_1 _07452_ (.A(net3212),
    .B(net856),
    .X(_00294_));
 sky130_fd_sc_hd__nor2_1 _07453_ (.A(_01769_),
    .B(net893),
    .Y(_00295_));
 sky130_fd_sc_hd__and2_1 _07454_ (.A(net3236),
    .B(net856),
    .X(_00296_));
 sky130_fd_sc_hd__and2_1 _07455_ (.A(net3116),
    .B(net856),
    .X(_00297_));
 sky130_fd_sc_hd__and2_1 _07456_ (.A(net3240),
    .B(net858),
    .X(_00298_));
 sky130_fd_sc_hd__nor2_1 _07457_ (.A(net3204),
    .B(net890),
    .Y(_00299_));
 sky130_fd_sc_hd__nor2_1 _07458_ (.A(net1173),
    .B(net890),
    .Y(_00300_));
 sky130_fd_sc_hd__nor2_1 _07459_ (.A(net3201),
    .B(net890),
    .Y(_00301_));
 sky130_fd_sc_hd__nor2_1 _07460_ (.A(net2951),
    .B(net890),
    .Y(_00302_));
 sky130_fd_sc_hd__and2_1 _07461_ (.A(net3086),
    .B(net856),
    .X(_00303_));
 sky130_fd_sc_hd__and2_1 _07462_ (.A(net1132),
    .B(net857),
    .X(_00304_));
 sky130_fd_sc_hd__and2_1 _07463_ (.A(net1168),
    .B(net857),
    .X(_00305_));
 sky130_fd_sc_hd__and2_1 _07464_ (.A(net875),
    .B(net944),
    .X(_00306_));
 sky130_fd_sc_hd__and2_1 _07465_ (.A(net876),
    .B(net924),
    .X(_00307_));
 sky130_fd_sc_hd__and2_1 _07466_ (.A(net876),
    .B(net932),
    .X(_00308_));
 sky130_fd_sc_hd__and2_1 _07467_ (.A(net876),
    .B(net922),
    .X(_00309_));
 sky130_fd_sc_hd__and2_1 _07468_ (.A(net857),
    .B(net1006),
    .X(_00310_));
 sky130_fd_sc_hd__and2_1 _07469_ (.A(net1040),
    .B(net856),
    .X(_00311_));
 sky130_fd_sc_hd__and2_1 _07470_ (.A(net1216),
    .B(net856),
    .X(_00312_));
 sky130_fd_sc_hd__and2_1 _07471_ (.A(net1152),
    .B(net861),
    .X(_00313_));
 sky130_fd_sc_hd__and2_1 _07472_ (.A(net1116),
    .B(net860),
    .X(_00314_));
 sky130_fd_sc_hd__and2_1 _07473_ (.A(net1138),
    .B(net861),
    .X(_00315_));
 sky130_fd_sc_hd__and2_1 _07474_ (.A(net1162),
    .B(net860),
    .X(_00316_));
 sky130_fd_sc_hd__and2_1 _07475_ (.A(net960),
    .B(net856),
    .X(_00317_));
 sky130_fd_sc_hd__or3_4 _07476_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(\ctrl.c2d_rf_waddr_W[3] ),
    .C(_01780_),
    .X(_02012_));
 sky130_fd_sc_hd__nor2_4 _07477_ (.A(_01821_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__mux2_1 _07478_ (.A0(net1880),
    .A1(net719),
    .S(net401),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _07479_ (.A0(net1790),
    .A1(net716),
    .S(net401),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _07480_ (.A0(net1412),
    .A1(net715),
    .S(net401),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _07481_ (.A0(net1922),
    .A1(net713),
    .S(net401),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _07482_ (.A0(net2322),
    .A1(net711),
    .S(net401),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _07483_ (.A0(net2008),
    .A1(net709),
    .S(net401),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _07484_ (.A0(net2426),
    .A1(net707),
    .S(net401),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _07485_ (.A0(net1988),
    .A1(net704),
    .S(net401),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _07486_ (.A0(net3709),
    .A1(net1180),
    .S(net401),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _07487_ (.A0(net2348),
    .A1(net701),
    .S(net401),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _07488_ (.A0(net1456),
    .A1(net699),
    .S(net401),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _07489_ (.A0(net2746),
    .A1(net696),
    .S(net401),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _07490_ (.A0(net2422),
    .A1(net695),
    .S(net401),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _07491_ (.A0(net2622),
    .A1(net692),
    .S(net401),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _07492_ (.A0(net2706),
    .A1(net691),
    .S(net401),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _07493_ (.A0(net1752),
    .A1(net689),
    .S(net401),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _07494_ (.A0(net1978),
    .A1(net687),
    .S(net402),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _07495_ (.A0(net2588),
    .A1(net685),
    .S(net402),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _07496_ (.A0(net2064),
    .A1(net683),
    .S(net402),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _07497_ (.A0(net2642),
    .A1(net680),
    .S(net402),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _07498_ (.A0(net1836),
    .A1(net678),
    .S(net402),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _07499_ (.A0(net2758),
    .A1(net675),
    .S(net402),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _07500_ (.A0(net2566),
    .A1(net674),
    .S(net402),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _07501_ (.A0(net2938),
    .A1(net672),
    .S(net402),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _07502_ (.A0(net2578),
    .A1(net668),
    .S(net402),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _07503_ (.A0(net2370),
    .A1(net666),
    .S(net402),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _07504_ (.A0(net1902),
    .A1(net664),
    .S(net402),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _07505_ (.A0(net1654),
    .A1(net662),
    .S(net402),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _07506_ (.A0(net2520),
    .A1(net660),
    .S(net402),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _07507_ (.A0(net2134),
    .A1(net658),
    .S(net402),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _07508_ (.A0(net2802),
    .A1(net656),
    .S(net402),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _07509_ (.A0(net2816),
    .A1(net654),
    .S(net402),
    .X(_00349_));
 sky130_fd_sc_hd__and3_2 _07510_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(_01779_),
    .C(\ctrl.c2d_rf_waddr_W[4] ),
    .X(_02014_));
 sky130_fd_sc_hd__or3_2 _07511_ (.A(_01778_),
    .B(\ctrl.c2d_rf_waddr_W[3] ),
    .C(_01780_),
    .X(_02015_));
 sky130_fd_sc_hd__nor2_4 _07512_ (.A(_01823_),
    .B(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__mux2_1 _07513_ (.A0(net1286),
    .A1(net719),
    .S(net439),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _07514_ (.A0(net1898),
    .A1(net3711),
    .S(net439),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _07515_ (.A0(net3000),
    .A1(net715),
    .S(net439),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _07516_ (.A0(net1254),
    .A1(net713),
    .S(net439),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _07517_ (.A0(net1646),
    .A1(net711),
    .S(net439),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _07518_ (.A0(net2574),
    .A1(net709),
    .S(net439),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _07519_ (.A0(net3188),
    .A1(net707),
    .S(net439),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _07520_ (.A0(net2128),
    .A1(net705),
    .S(net439),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _07521_ (.A0(net2722),
    .A1(net702),
    .S(net439),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _07522_ (.A0(net2824),
    .A1(net701),
    .S(net439),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _07523_ (.A0(net1794),
    .A1(net699),
    .S(net439),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _07524_ (.A0(net2540),
    .A1(net696),
    .S(net439),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _07525_ (.A0(net1450),
    .A1(net3717),
    .S(net439),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _07526_ (.A0(net1960),
    .A1(net692),
    .S(net439),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(net1596),
    .A1(net691),
    .S(net439),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _07528_ (.A0(net1500),
    .A1(net689),
    .S(net439),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _07529_ (.A0(net2010),
    .A1(net687),
    .S(net440),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _07530_ (.A0(net3700),
    .A1(net1064),
    .S(net440),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _07531_ (.A0(net1200),
    .A1(net683),
    .S(net440),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _07532_ (.A0(net1312),
    .A1(net681),
    .S(net440),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _07533_ (.A0(net1410),
    .A1(net679),
    .S(net440),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _07534_ (.A0(net1284),
    .A1(net676),
    .S(net440),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _07535_ (.A0(net1586),
    .A1(net3714),
    .S(net440),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _07536_ (.A0(net1540),
    .A1(net672),
    .S(net440),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _07537_ (.A0(net1362),
    .A1(net670),
    .S(net440),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _07538_ (.A0(net1372),
    .A1(net667),
    .S(net440),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _07539_ (.A0(net2494),
    .A1(net664),
    .S(net440),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _07540_ (.A0(net1528),
    .A1(net663),
    .S(net440),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _07541_ (.A0(net1388),
    .A1(net660),
    .S(net440),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _07542_ (.A0(net1720),
    .A1(net659),
    .S(net440),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _07543_ (.A0(net1252),
    .A1(net656),
    .S(net440),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _07544_ (.A0(net2130),
    .A1(net655),
    .S(net440),
    .X(_00381_));
 sky130_fd_sc_hd__and2_1 _07545_ (.A(net847),
    .B(net1068),
    .X(_00382_));
 sky130_fd_sc_hd__and2_1 _07546_ (.A(net847),
    .B(net908),
    .X(_00383_));
 sky130_fd_sc_hd__and2_1 _07547_ (.A(net847),
    .B(net1084),
    .X(_00384_));
 sky130_fd_sc_hd__and2_1 _07548_ (.A(net847),
    .B(net1106),
    .X(_00385_));
 sky130_fd_sc_hd__and2_1 _07549_ (.A(net847),
    .B(net1128),
    .X(_00386_));
 sky130_fd_sc_hd__and2_1 _07550_ (.A(net847),
    .B(net1110),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _07551_ (.A(net847),
    .B(net1070),
    .X(_00388_));
 sky130_fd_sc_hd__and2_1 _07552_ (.A(net848),
    .B(net986),
    .X(_00389_));
 sky130_fd_sc_hd__and2_1 _07553_ (.A(net848),
    .B(net1046),
    .X(_00390_));
 sky130_fd_sc_hd__and2_1 _07554_ (.A(net847),
    .B(net1026),
    .X(_00391_));
 sky130_fd_sc_hd__and2_1 _07555_ (.A(net848),
    .B(net3206),
    .X(_00392_));
 sky130_fd_sc_hd__and2_1 _07556_ (.A(net848),
    .B(net1030),
    .X(_00393_));
 sky130_fd_sc_hd__and2_1 _07557_ (.A(net848),
    .B(net1024),
    .X(_00394_));
 sky130_fd_sc_hd__and2_1 _07558_ (.A(net848),
    .B(net1044),
    .X(_00395_));
 sky130_fd_sc_hd__and2_1 _07559_ (.A(net848),
    .B(net1038),
    .X(_00396_));
 sky130_fd_sc_hd__and2_1 _07560_ (.A(net848),
    .B(net1020),
    .X(_00397_));
 sky130_fd_sc_hd__and2_1 _07561_ (.A(net863),
    .B(net1072),
    .X(_00398_));
 sky130_fd_sc_hd__and2_1 _07562_ (.A(net863),
    .B(net1014),
    .X(_00399_));
 sky130_fd_sc_hd__and2_1 _07563_ (.A(net863),
    .B(net1086),
    .X(_00400_));
 sky130_fd_sc_hd__and2_1 _07564_ (.A(net863),
    .B(net1034),
    .X(_00401_));
 sky130_fd_sc_hd__and2_1 _07565_ (.A(net863),
    .B(net1076),
    .X(_00402_));
 sky130_fd_sc_hd__and2_1 _07566_ (.A(net863),
    .B(net1104),
    .X(_00403_));
 sky130_fd_sc_hd__and2_1 _07567_ (.A(net863),
    .B(net1088),
    .X(_00404_));
 sky130_fd_sc_hd__and2_1 _07568_ (.A(net863),
    .B(net1050),
    .X(_00405_));
 sky130_fd_sc_hd__and2_1 _07569_ (.A(net863),
    .B(net1056),
    .X(_00406_));
 sky130_fd_sc_hd__and2_1 _07570_ (.A(net864),
    .B(net1062),
    .X(_00407_));
 sky130_fd_sc_hd__and2_1 _07571_ (.A(net863),
    .B(net3288),
    .X(_00408_));
 sky130_fd_sc_hd__and2_1 _07572_ (.A(net863),
    .B(net3425),
    .X(_00409_));
 sky130_fd_sc_hd__and2_1 _07573_ (.A(net865),
    .B(net3442),
    .X(_00410_));
 sky130_fd_sc_hd__and2_1 _07574_ (.A(net865),
    .B(net3244),
    .X(_00411_));
 sky130_fd_sc_hd__and2_1 _07575_ (.A(net865),
    .B(net3270),
    .X(_00412_));
 sky130_fd_sc_hd__and2_1 _07576_ (.A(net865),
    .B(net3308),
    .X(_00413_));
 sky130_fd_sc_hd__nand2_4 _07577_ (.A(_01829_),
    .B(_02014_),
    .Y(_02017_));
 sky130_fd_sc_hd__mux2_1 _07578_ (.A0(net719),
    .A1(net2078),
    .S(net399),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _07579_ (.A0(net716),
    .A1(net1392),
    .S(net399),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _07580_ (.A0(net715),
    .A1(net2532),
    .S(net399),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _07581_ (.A0(net713),
    .A1(net2634),
    .S(net399),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _07582_ (.A0(net711),
    .A1(net2380),
    .S(net399),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _07583_ (.A0(net709),
    .A1(net2590),
    .S(net399),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _07584_ (.A0(net707),
    .A1(net2988),
    .S(net399),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _07585_ (.A0(\dpath.RF.wdata[7] ),
    .A1(net1696),
    .S(net399),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _07586_ (.A0(net702),
    .A1(net1390),
    .S(net399),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _07587_ (.A0(net701),
    .A1(net1472),
    .S(net399),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _07588_ (.A0(net699),
    .A1(net1944),
    .S(net399),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _07589_ (.A0(net696),
    .A1(net2560),
    .S(net399),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _07590_ (.A0(net3717),
    .A1(net2828),
    .S(net399),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _07591_ (.A0(net692),
    .A1(net2038),
    .S(net399),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _07592_ (.A0(net691),
    .A1(net2964),
    .S(net399),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _07593_ (.A0(net689),
    .A1(net2362),
    .S(net399),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _07594_ (.A0(net687),
    .A1(net1906),
    .S(net400),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _07595_ (.A0(net685),
    .A1(net2098),
    .S(net400),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _07596_ (.A0(\dpath.RF.wdata[18] ),
    .A1(net2800),
    .S(net400),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _07597_ (.A0(net998),
    .A1(net3713),
    .S(net400),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _07598_ (.A0(net678),
    .A1(net2318),
    .S(net400),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _07599_ (.A0(net676),
    .A1(net2598),
    .S(net400),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _07600_ (.A0(net674),
    .A1(net3060),
    .S(net400),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _07601_ (.A0(net672),
    .A1(net2188),
    .S(net400),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _07602_ (.A0(net668),
    .A1(net3100),
    .S(net400),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _07603_ (.A0(net666),
    .A1(net2352),
    .S(net400),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _07604_ (.A0(net664),
    .A1(net2516),
    .S(net400),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _07605_ (.A0(net663),
    .A1(net2492),
    .S(net400),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _07606_ (.A0(net660),
    .A1(net1730),
    .S(net400),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _07607_ (.A0(net659),
    .A1(net3008),
    .S(net400),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _07608_ (.A0(net656),
    .A1(net1718),
    .S(net400),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _07609_ (.A0(net655),
    .A1(net2360),
    .S(net400),
    .X(_00445_));
 sky130_fd_sc_hd__nor2_4 _07610_ (.A(_01830_),
    .B(_02012_),
    .Y(_02018_));
 sky130_fd_sc_hd__mux2_1 _07611_ (.A0(net2924),
    .A1(net719),
    .S(net397),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _07612_ (.A0(net2980),
    .A1(net716),
    .S(net397),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _07613_ (.A0(net1222),
    .A1(net715),
    .S(net397),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _07614_ (.A0(net2726),
    .A1(net713),
    .S(net397),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _07615_ (.A0(net2412),
    .A1(net711),
    .S(net397),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _07616_ (.A0(net2886),
    .A1(net709),
    .S(net397),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _07617_ (.A0(net1808),
    .A1(net707),
    .S(net397),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _07618_ (.A0(net2262),
    .A1(net704),
    .S(net397),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _07619_ (.A0(net1628),
    .A1(net702),
    .S(net397),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _07620_ (.A0(net2286),
    .A1(net701),
    .S(net397),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _07621_ (.A0(net1726),
    .A1(net699),
    .S(net397),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _07622_ (.A0(net1868),
    .A1(net696),
    .S(net397),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _07623_ (.A0(net2714),
    .A1(net695),
    .S(net397),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _07624_ (.A0(net2730),
    .A1(net692),
    .S(net397),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _07625_ (.A0(net2820),
    .A1(net691),
    .S(net397),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _07626_ (.A0(net1496),
    .A1(net689),
    .S(net397),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _07627_ (.A0(net1440),
    .A1(net687),
    .S(net398),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _07628_ (.A0(net1956),
    .A1(net685),
    .S(net398),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _07629_ (.A0(net2602),
    .A1(net683),
    .S(net398),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _07630_ (.A0(net2328),
    .A1(net680),
    .S(net398),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _07631_ (.A0(net1428),
    .A1(net678),
    .S(net398),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _07632_ (.A0(net1976),
    .A1(net675),
    .S(net398),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _07633_ (.A0(net1594),
    .A1(net674),
    .S(net398),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _07634_ (.A0(net2314),
    .A1(net672),
    .S(net398),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(net2190),
    .A1(net668),
    .S(net398),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _07636_ (.A0(net1462),
    .A1(net666),
    .S(net398),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _07637_ (.A0(net1328),
    .A1(net664),
    .S(net398),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _07638_ (.A0(net1798),
    .A1(net662),
    .S(net398),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _07639_ (.A0(net1562),
    .A1(net660),
    .S(net398),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _07640_ (.A0(net1692),
    .A1(net658),
    .S(net398),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(net2336),
    .A1(net656),
    .S(net398),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _07642_ (.A0(net2686),
    .A1(net654),
    .S(net398),
    .X(_00477_));
 sky130_fd_sc_hd__or4b_4 _07643_ (.A(\ctrl.c2d_rf_waddr_W[0] ),
    .B(\ctrl.c2d_rf_waddr_W[1] ),
    .C(_01818_),
    .D_N(_01832_),
    .X(_02019_));
 sky130_fd_sc_hd__nor2_4 _07644_ (.A(_02015_),
    .B(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__mux2_1 _07645_ (.A0(net1514),
    .A1(net719),
    .S(net437),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _07646_ (.A0(net1404),
    .A1(net716),
    .S(net437),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _07647_ (.A0(net3098),
    .A1(net715),
    .S(net437),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _07648_ (.A0(net1318),
    .A1(net713),
    .S(net437),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _07649_ (.A0(net2076),
    .A1(net711),
    .S(net437),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _07650_ (.A0(net1398),
    .A1(net709),
    .S(net437),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _07651_ (.A0(net2454),
    .A1(net707),
    .S(net437),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _07652_ (.A0(net2934),
    .A1(\dpath.RF.wdata[7] ),
    .S(net437),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _07653_ (.A0(net1274),
    .A1(net703),
    .S(net437),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _07654_ (.A0(net2056),
    .A1(net701),
    .S(net437),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _07655_ (.A0(net1716),
    .A1(net699),
    .S(net437),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _07656_ (.A0(net1888),
    .A1(net696),
    .S(net437),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _07657_ (.A0(net1506),
    .A1(net695),
    .S(net437),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _07658_ (.A0(net2168),
    .A1(net692),
    .S(net437),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _07659_ (.A0(net1694),
    .A1(net691),
    .S(net437),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _07660_ (.A0(net1652),
    .A1(net689),
    .S(net437),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _07661_ (.A0(net2716),
    .A1(net687),
    .S(net438),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _07662_ (.A0(net2160),
    .A1(net1064),
    .S(net438),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _07663_ (.A0(net1568),
    .A1(\dpath.RF.wdata[18] ),
    .S(net438),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _07664_ (.A0(net2106),
    .A1(net680),
    .S(net438),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _07665_ (.A0(net1700),
    .A1(net678),
    .S(net438),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _07666_ (.A0(net1874),
    .A1(net676),
    .S(net438),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _07667_ (.A0(net1488),
    .A1(net674),
    .S(net438),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _07668_ (.A0(net2146),
    .A1(net672),
    .S(net438),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _07669_ (.A0(net1320),
    .A1(net668),
    .S(net438),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _07670_ (.A0(net2206),
    .A1(net666),
    .S(net438),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _07671_ (.A0(net2732),
    .A1(net3659),
    .S(net438),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _07672_ (.A0(net2756),
    .A1(net663),
    .S(net438),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _07673_ (.A0(net1494),
    .A1(net660),
    .S(net438),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _07674_ (.A0(net1708),
    .A1(\dpath.RF.wdata[29] ),
    .S(net438),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _07675_ (.A0(net2324),
    .A1(net656),
    .S(net438),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _07676_ (.A0(net2890),
    .A1(net655),
    .S(net438),
    .X(_00509_));
 sky130_fd_sc_hd__nor2_4 _07677_ (.A(_01830_),
    .B(_01832_),
    .Y(_02021_));
 sky130_fd_sc_hd__mux2_1 _07678_ (.A0(net1424),
    .A1(net718),
    .S(net395),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _07679_ (.A0(net1638),
    .A1(net717),
    .S(net395),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _07680_ (.A0(net1196),
    .A1(net714),
    .S(net395),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _07681_ (.A0(net1298),
    .A1(net712),
    .S(net395),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _07682_ (.A0(net2176),
    .A1(net710),
    .S(net395),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _07683_ (.A0(net2482),
    .A1(net708),
    .S(net395),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _07684_ (.A0(net1228),
    .A1(net706),
    .S(net395),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _07685_ (.A0(net1240),
    .A1(net705),
    .S(net395),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _07686_ (.A0(net2026),
    .A1(net702),
    .S(net395),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _07687_ (.A0(net2586),
    .A1(net700),
    .S(net395),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _07688_ (.A0(net1400),
    .A1(net698),
    .S(net395),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _07689_ (.A0(net1712),
    .A1(net697),
    .S(net395),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _07690_ (.A0(net1260),
    .A1(net694),
    .S(net395),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _07691_ (.A0(net2394),
    .A1(net693),
    .S(net395),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _07692_ (.A0(net2180),
    .A1(net690),
    .S(net395),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _07693_ (.A0(net2344),
    .A1(net688),
    .S(net395),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _07694_ (.A0(net2020),
    .A1(net686),
    .S(net396),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _07695_ (.A0(net1532),
    .A1(net684),
    .S(net396),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _07696_ (.A0(net1966),
    .A1(net682),
    .S(net396),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _07697_ (.A0(net1432),
    .A1(net681),
    .S(net396),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _07698_ (.A0(net2766),
    .A1(net677),
    .S(net396),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _07699_ (.A0(net2544),
    .A1(net675),
    .S(net396),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _07700_ (.A0(net1454),
    .A1(net673),
    .S(net396),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _07701_ (.A0(net1230),
    .A1(net671),
    .S(net396),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _07702_ (.A0(net1192),
    .A1(net669),
    .S(net396),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _07703_ (.A0(net1522),
    .A1(net666),
    .S(net396),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _07704_ (.A0(net1856),
    .A1(net665),
    .S(net396),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _07705_ (.A0(net2778),
    .A1(net662),
    .S(net396),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _07706_ (.A0(net1212),
    .A1(net661),
    .S(net396),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _07707_ (.A0(net1426),
    .A1(net658),
    .S(net396),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _07708_ (.A0(net2124),
    .A1(net657),
    .S(net396),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _07709_ (.A0(net2114),
    .A1(net654),
    .S(net396),
    .X(_00541_));
 sky130_fd_sc_hd__and3b_4 _07710_ (.A_N(_02019_),
    .B(_01779_),
    .C(_01778_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _07711_ (.A0(net2158),
    .A1(net719),
    .S(net435),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _07712_ (.A0(net3050),
    .A1(net716),
    .S(net435),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _07713_ (.A0(net1420),
    .A1(net715),
    .S(net435),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _07714_ (.A0(net1490),
    .A1(net713),
    .S(net435),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _07715_ (.A0(net1498),
    .A1(net711),
    .S(net435),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _07716_ (.A0(net1310),
    .A1(net709),
    .S(net435),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _07717_ (.A0(net1232),
    .A1(net707),
    .S(net435),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _07718_ (.A0(net1746),
    .A1(net704),
    .S(net435),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _07719_ (.A0(net1356),
    .A1(net702),
    .S(net435),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _07720_ (.A0(net1394),
    .A1(net701),
    .S(net435),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _07721_ (.A0(net1214),
    .A1(net699),
    .S(net435),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _07722_ (.A0(net1526),
    .A1(net696),
    .S(net435),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _07723_ (.A0(net2004),
    .A1(net695),
    .S(net435),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _07724_ (.A0(net1884),
    .A1(net692),
    .S(net435),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _07725_ (.A0(net2242),
    .A1(net691),
    .S(net435),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _07726_ (.A0(net1358),
    .A1(net689),
    .S(net435),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _07727_ (.A0(net1434),
    .A1(net687),
    .S(net436),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _07728_ (.A0(net2570),
    .A1(net685),
    .S(net436),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _07729_ (.A0(net2514),
    .A1(net683),
    .S(net436),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _07730_ (.A0(net2448),
    .A1(net680),
    .S(net436),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _07731_ (.A0(net1302),
    .A1(net677),
    .S(net436),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _07732_ (.A0(net1278),
    .A1(net675),
    .S(net436),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _07733_ (.A0(net1826),
    .A1(net674),
    .S(net436),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _07734_ (.A0(net2264),
    .A1(net672),
    .S(net436),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _07735_ (.A0(net2456),
    .A1(net668),
    .S(net436),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _07736_ (.A0(net2350),
    .A1(net666),
    .S(net436),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _07737_ (.A0(net3038),
    .A1(net664),
    .S(net436),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _07738_ (.A0(net1630),
    .A1(net662),
    .S(net436),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _07739_ (.A0(net1990),
    .A1(net660),
    .S(net436),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _07740_ (.A0(net1524),
    .A1(net659),
    .S(net436),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _07741_ (.A0(net1552),
    .A1(net656),
    .S(net436),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _07742_ (.A0(net2358),
    .A1(net654),
    .S(net436),
    .X(_00573_));
 sky130_fd_sc_hd__and3_2 _07743_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(\ctrl.c2d_rf_waddr_W[3] ),
    .C(_01780_),
    .X(_02023_));
 sky130_fd_sc_hd__or3_2 _07744_ (.A(_01778_),
    .B(_01779_),
    .C(\ctrl.c2d_rf_waddr_W[4] ),
    .X(_02024_));
 sky130_fd_sc_hd__nand2_4 _07745_ (.A(_01820_),
    .B(_02023_),
    .Y(_02025_));
 sky130_fd_sc_hd__mux2_1 _07746_ (.A0(net718),
    .A1(net3018),
    .S(net393),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _07747_ (.A0(net717),
    .A1(net3036),
    .S(net393),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _07748_ (.A0(net714),
    .A1(net2254),
    .S(net393),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _07749_ (.A0(net712),
    .A1(net2104),
    .S(net393),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _07750_ (.A0(net710),
    .A1(net3032),
    .S(net393),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _07751_ (.A0(net708),
    .A1(net2908),
    .S(net393),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _07752_ (.A0(net707),
    .A1(net2608),
    .S(net393),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _07753_ (.A0(net704),
    .A1(net2880),
    .S(net393),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _07754_ (.A0(net703),
    .A1(net1352),
    .S(net393),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _07755_ (.A0(net700),
    .A1(net2016),
    .S(net393),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _07756_ (.A0(net698),
    .A1(net3034),
    .S(net393),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _07757_ (.A0(net697),
    .A1(net2604),
    .S(net393),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _07758_ (.A0(net694),
    .A1(net2724),
    .S(net393),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _07759_ (.A0(net693),
    .A1(net2488),
    .S(net393),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _07760_ (.A0(net690),
    .A1(net2266),
    .S(net393),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _07761_ (.A0(net688),
    .A1(net2678),
    .S(net393),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _07762_ (.A0(net686),
    .A1(net2946),
    .S(net394),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _07763_ (.A0(net684),
    .A1(net2268),
    .S(net394),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _07764_ (.A0(net682),
    .A1(net3014),
    .S(net394),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _07765_ (.A0(net680),
    .A1(net2108),
    .S(net394),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _07766_ (.A0(net677),
    .A1(net3138),
    .S(net394),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _07767_ (.A0(net675),
    .A1(net2858),
    .S(net394),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _07768_ (.A0(net673),
    .A1(net2936),
    .S(net394),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _07769_ (.A0(net671),
    .A1(net2882),
    .S(net394),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _07770_ (.A0(net669),
    .A1(net2870),
    .S(net394),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _07771_ (.A0(net666),
    .A1(net2872),
    .S(net394),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _07772_ (.A0(net665),
    .A1(net2676),
    .S(net394),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _07773_ (.A0(net662),
    .A1(net2862),
    .S(net394),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _07774_ (.A0(net661),
    .A1(net2430),
    .S(net394),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _07775_ (.A0(net658),
    .A1(net2240),
    .S(net394),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _07776_ (.A0(net657),
    .A1(net2024),
    .S(net394),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _07777_ (.A0(net654),
    .A1(net2174),
    .S(net394),
    .X(_00605_));
 sky130_fd_sc_hd__nor2_4 _07778_ (.A(_01823_),
    .B(_02012_),
    .Y(_02026_));
 sky130_fd_sc_hd__mux2_1 _07779_ (.A0(net1486),
    .A1(net719),
    .S(net433),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _07780_ (.A0(net1986),
    .A1(net716),
    .S(net433),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _07781_ (.A0(net2220),
    .A1(net715),
    .S(net433),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _07782_ (.A0(net1276),
    .A1(net713),
    .S(net433),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _07783_ (.A0(net1674),
    .A1(net711),
    .S(net433),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _07784_ (.A0(net2186),
    .A1(net709),
    .S(net433),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _07785_ (.A0(net2630),
    .A1(net707),
    .S(net433),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _07786_ (.A0(net1336),
    .A1(net704),
    .S(net433),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _07787_ (.A0(net1304),
    .A1(net702),
    .S(net433),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _07788_ (.A0(net1820),
    .A1(net701),
    .S(net433),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _07789_ (.A0(net1854),
    .A1(net699),
    .S(net433),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _07790_ (.A0(net1676),
    .A1(net696),
    .S(net433),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _07791_ (.A0(net2760),
    .A1(net695),
    .S(net433),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _07792_ (.A0(net1864),
    .A1(net692),
    .S(net433),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _07793_ (.A0(net2728),
    .A1(net691),
    .S(net433),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _07794_ (.A0(net1642),
    .A1(net689),
    .S(net433),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _07795_ (.A0(net2310),
    .A1(net687),
    .S(net434),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _07796_ (.A0(net1872),
    .A1(net685),
    .S(net434),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _07797_ (.A0(net1478),
    .A1(net683),
    .S(net434),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _07798_ (.A0(net1370),
    .A1(net680),
    .S(net434),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _07799_ (.A0(net1538),
    .A1(net678),
    .S(net434),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _07800_ (.A0(net2022),
    .A1(net675),
    .S(net434),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _07801_ (.A0(net1396),
    .A1(net674),
    .S(net434),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _07802_ (.A0(net1736),
    .A1(net672),
    .S(net434),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _07803_ (.A0(net1792),
    .A1(net668),
    .S(net434),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _07804_ (.A0(net1442),
    .A1(net666),
    .S(net434),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _07805_ (.A0(net3108),
    .A1(net664),
    .S(net434),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _07806_ (.A0(net1204),
    .A1(net662),
    .S(net434),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _07807_ (.A0(net1974),
    .A1(net660),
    .S(net434),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _07808_ (.A0(net1384),
    .A1(net659),
    .S(net434),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _07809_ (.A0(net1368),
    .A1(net656),
    .S(net434),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _07810_ (.A0(net1780),
    .A1(net654),
    .S(net434),
    .X(_00637_));
 sky130_fd_sc_hd__nor2_4 _07811_ (.A(net404),
    .B(_01955_),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_1 _07812_ (.A(net404),
    .B(_01955_),
    .X(_02028_));
 sky130_fd_sc_hd__mux4_1 _07813_ (.A0(\dpath.RF.R[0][2] ),
    .A1(\dpath.RF.R[1][2] ),
    .A2(\dpath.RF.R[2][2] ),
    .A3(\dpath.RF.R[3][2] ),
    .S0(net563),
    .S1(net543),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _07814_ (.A0(\dpath.RF.R[6][2] ),
    .A1(\dpath.RF.R[7][2] ),
    .S(net564),
    .X(_02030_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(net545),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__mux2_1 _07816_ (.A0(\dpath.RF.R[4][2] ),
    .A1(\dpath.RF.R[5][2] ),
    .S(net564),
    .X(_02032_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(_01770_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__o21ai_1 _07818_ (.A1(net531),
    .A2(_02029_),
    .B1(net506),
    .Y(_02034_));
 sky130_fd_sc_hd__a31o_1 _07819_ (.A1(net531),
    .A2(_02031_),
    .A3(_02033_),
    .B1(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__mux4_1 _07820_ (.A0(\dpath.RF.R[12][2] ),
    .A1(\dpath.RF.R[13][2] ),
    .A2(\dpath.RF.R[14][2] ),
    .A3(\dpath.RF.R[15][2] ),
    .S0(net562),
    .S1(net543),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _07821_ (.A0(\dpath.RF.R[8][2] ),
    .A1(\dpath.RF.R[9][2] ),
    .S(net565),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _07822_ (.A0(\dpath.RF.R[10][2] ),
    .A1(\dpath.RF.R[11][2] ),
    .S(net565),
    .X(_02038_));
 sky130_fd_sc_hd__a21o_1 _07823_ (.A1(net544),
    .A2(_02038_),
    .B1(net532),
    .X(_02039_));
 sky130_fd_sc_hd__a21o_1 _07824_ (.A1(_01770_),
    .A2(_02037_),
    .B1(_02039_),
    .X(_02040_));
 sky130_fd_sc_hd__o211a_1 _07825_ (.A1(net511),
    .A2(_02036_),
    .B1(_02040_),
    .C1(net523),
    .X(_02041_));
 sky130_fd_sc_hd__nor2_1 _07826_ (.A(net518),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__mux4_1 _07827_ (.A0(\dpath.RF.R[16][2] ),
    .A1(\dpath.RF.R[17][2] ),
    .A2(\dpath.RF.R[18][2] ),
    .A3(\dpath.RF.R[19][2] ),
    .S0(net564),
    .S1(net545),
    .X(_02043_));
 sky130_fd_sc_hd__nor2_1 _07828_ (.A(net532),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__mux4_1 _07829_ (.A0(\dpath.RF.R[20][2] ),
    .A1(\dpath.RF.R[21][2] ),
    .A2(\dpath.RF.R[22][2] ),
    .A3(\dpath.RF.R[23][2] ),
    .S0(net562),
    .S1(net546),
    .X(_02045_));
 sky130_fd_sc_hd__nor2_1 _07830_ (.A(net511),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__mux4_1 _07831_ (.A0(\dpath.RF.R[28][2] ),
    .A1(\dpath.RF.R[29][2] ),
    .A2(\dpath.RF.R[30][2] ),
    .A3(\dpath.RF.R[31][2] ),
    .S0(net564),
    .S1(net545),
    .X(_02047_));
 sky130_fd_sc_hd__nor2_1 _07832_ (.A(net511),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__mux4_1 _07833_ (.A0(\dpath.RF.R[24][2] ),
    .A1(\dpath.RF.R[25][2] ),
    .A2(\dpath.RF.R[26][2] ),
    .A3(\dpath.RF.R[27][2] ),
    .S0(net563),
    .S1(net543),
    .X(_02049_));
 sky130_fd_sc_hd__o21ai_1 _07834_ (.A1(net531),
    .A2(_02049_),
    .B1(net523),
    .Y(_02050_));
 sky130_fd_sc_hd__o32a_1 _07835_ (.A1(net523),
    .A2(_02044_),
    .A3(_02046_),
    .B1(_02048_),
    .B2(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__a22o_1 _07836_ (.A1(_02035_),
    .A2(_02042_),
    .B1(_02051_),
    .B2(net518),
    .X(_02052_));
 sky130_fd_sc_hd__o31ai_2 _07837_ (.A1(\ctrl.inst_M[4] ),
    .A2(\ctrl.inst_M[5] ),
    .A3(_01796_),
    .B1(_01804_),
    .Y(_02053_));
 sky130_fd_sc_hd__xnor2_1 _07838_ (.A(\ctrl.d2c_inst[17] ),
    .B(\ctrl.inst_M[9] ),
    .Y(_02054_));
 sky130_fd_sc_hd__o2bb2a_1 _07839_ (.A1_N(_01758_),
    .A2_N(\ctrl.inst_M[7] ),
    .B1(\ctrl.inst_M[10] ),
    .B2(_01755_),
    .X(_02055_));
 sky130_fd_sc_hd__or3_1 _07840_ (.A(\ctrl.inst_M[9] ),
    .B(\ctrl.inst_M[10] ),
    .C(\ctrl.inst_M[11] ),
    .X(_02056_));
 sky130_fd_sc_hd__or3_1 _07841_ (.A(\ctrl.inst_M[7] ),
    .B(\ctrl.inst_M[8] ),
    .C(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__o221a_1 _07842_ (.A1(_01758_),
    .A2(\ctrl.inst_M[7] ),
    .B1(\ctrl.inst_M[11] ),
    .B2(_01754_),
    .C1(_02055_),
    .X(_02058_));
 sky130_fd_sc_hd__o2111a_1 _07843_ (.A1(\ctrl.d2c_inst[16] ),
    .A2(_01781_),
    .B1(_02054_),
    .C1(_02058_),
    .D1(\ctrl.val_M ),
    .X(_02059_));
 sky130_fd_sc_hd__o22a_1 _07844_ (.A1(\ctrl.d2c_inst[18] ),
    .A2(_01783_),
    .B1(_01784_),
    .B2(\ctrl.d2c_inst[19] ),
    .X(_02060_));
 sky130_fd_sc_hd__o2111a_1 _07845_ (.A1(_01757_),
    .A2(\ctrl.inst_M[8] ),
    .B1(_02057_),
    .C1(_02059_),
    .D1(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__nand3_1 _07846_ (.A(_01981_),
    .B(_02053_),
    .C(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__or4_1 _07847_ (.A(\ctrl.inst_X[28] ),
    .B(\ctrl.inst_X[27] ),
    .C(\ctrl.inst_X[30] ),
    .D(\ctrl.inst_X[29] ),
    .X(_02063_));
 sky130_fd_sc_hd__o41a_1 _07848_ (.A1(\ctrl.inst_X[31] ),
    .A2(\ctrl.inst_X[26] ),
    .A3(\ctrl.inst_X[25] ),
    .A4(_02063_),
    .B1(\ctrl.inst_X[5] ),
    .X(_02064_));
 sky130_fd_sc_hd__and4b_1 _07849_ (.A_N(_02064_),
    .B(_01959_),
    .C(_01839_),
    .D(\ctrl.inst_X[4] ),
    .X(_02065_));
 sky130_fd_sc_hd__and4_1 _07850_ (.A(\ctrl.inst_X[1] ),
    .B(\ctrl.inst_X[0] ),
    .C(\ctrl.inst_X[3] ),
    .D(\ctrl.inst_X[2] ),
    .X(_02066_));
 sky130_fd_sc_hd__a21oi_4 _07851_ (.A1(_01838_),
    .A2(_02066_),
    .B1(_02065_),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _07852_ (.A(net3207),
    .B(net3209),
    .Y(_02068_));
 sky130_fd_sc_hd__or4bb_1 _07853_ (.A(\ctrl.inst_X[12] ),
    .B(\ctrl.inst_X[14] ),
    .C_N(\ctrl.inst_X[13] ),
    .D_N(\ctrl.inst_X[6] ),
    .X(_02069_));
 sky130_fd_sc_hd__nor3_2 _07854_ (.A(_01837_),
    .B(_02068_),
    .C(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__or3_4 _07855_ (.A(_01837_),
    .B(_02068_),
    .C(_02069_),
    .X(_02071_));
 sky130_fd_sc_hd__nand2_1 _07856_ (.A(\ctrl.inst_X[25] ),
    .B(_01839_),
    .Y(_02072_));
 sky130_fd_sc_hd__or4_1 _07857_ (.A(\ctrl.inst_X[31] ),
    .B(\ctrl.inst_X[26] ),
    .C(_02068_),
    .D(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__o311a_1 _07858_ (.A1(_01960_),
    .A2(_02063_),
    .A3(_02073_),
    .B1(net484),
    .C1(_02067_),
    .X(_02074_));
 sky130_fd_sc_hd__inv_2 _07859_ (.A(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__o211a_2 _07860_ (.A1(\ctrl.inst_X[9] ),
    .A2(_01963_),
    .B1(_02075_),
    .C1(_01962_),
    .X(_02076_));
 sky130_fd_sc_hd__nor2_1 _07861_ (.A(\ctrl.d2c_inst[19] ),
    .B(\ctrl.d2c_inst[18] ),
    .Y(_02077_));
 sky130_fd_sc_hd__and4_4 _07862_ (.A(_01756_),
    .B(_01757_),
    .C(_01758_),
    .D(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__nand3_1 _07863_ (.A(\ctrl.inst_W[5] ),
    .B(\ctrl.inst_W[4] ),
    .C(\ctrl.inst_W[6] ),
    .Y(_02079_));
 sky130_fd_sc_hd__or3_1 _07864_ (.A(\ctrl.inst_W[5] ),
    .B(\ctrl.inst_W[4] ),
    .C(\ctrl.inst_W[6] ),
    .X(_02080_));
 sky130_fd_sc_hd__a211o_1 _07865_ (.A1(_02079_),
    .A2(_02080_),
    .B1(\ctrl.inst_W[14] ),
    .C1(_01775_),
    .X(_02081_));
 sky130_fd_sc_hd__or4_1 _07866_ (.A(\ctrl.inst_W[28] ),
    .B(\ctrl.inst_W[30] ),
    .C(\ctrl.inst_W[29] ),
    .D(\ctrl.inst_W[31] ),
    .X(_02082_));
 sky130_fd_sc_hd__o31a_1 _07867_ (.A1(\ctrl.inst_W[26] ),
    .A2(\ctrl.inst_W[27] ),
    .A3(_02082_),
    .B1(\ctrl.inst_W[5] ),
    .X(_02083_));
 sky130_fd_sc_hd__or3b_1 _07868_ (.A(\ctrl.inst_W[14] ),
    .B(\ctrl.inst_W[13] ),
    .C_N(\ctrl.inst_W[4] ),
    .X(_02084_));
 sky130_fd_sc_hd__o31a_1 _07869_ (.A1(\ctrl.inst_W[6] ),
    .A2(_02083_),
    .A3(_02084_),
    .B1(_02081_),
    .X(_02085_));
 sky130_fd_sc_hd__o32a_1 _07870_ (.A1(\ctrl.inst_W[12] ),
    .A2(_01812_),
    .A3(_02085_),
    .B1(_01811_),
    .B2(_01774_),
    .X(_02086_));
 sky130_fd_sc_hd__a22o_1 _07871_ (.A1(_01757_),
    .A2(\ctrl.c2d_rf_waddr_W[1] ),
    .B1(_01778_),
    .B2(\ctrl.d2c_inst[17] ),
    .X(_02087_));
 sky130_fd_sc_hd__a221o_1 _07872_ (.A1(_01756_),
    .A2(\ctrl.c2d_rf_waddr_W[2] ),
    .B1(_01780_),
    .B2(\ctrl.d2c_inst[19] ),
    .C1(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__a22o_1 _07873_ (.A1(\ctrl.d2c_inst[16] ),
    .A2(_01777_),
    .B1(\ctrl.c2d_rf_waddr_W[3] ),
    .B2(_01755_),
    .X(_02089_));
 sky130_fd_sc_hd__a2111o_1 _07874_ (.A1(\ctrl.d2c_inst[18] ),
    .A2(_01779_),
    .B1(_02088_),
    .C1(_02089_),
    .D1(_01773_),
    .X(_02090_));
 sky130_fd_sc_hd__and3b_1 _07875_ (.A_N(_01832_),
    .B(_01777_),
    .C(_01776_),
    .X(_02091_));
 sky130_fd_sc_hd__a22o_1 _07876_ (.A1(\ctrl.d2c_inst[15] ),
    .A2(_01776_),
    .B1(\ctrl.c2d_rf_waddr_W[4] ),
    .B2(_01754_),
    .X(_02092_));
 sky130_fd_sc_hd__a211o_1 _07877_ (.A1(_01758_),
    .A2(\ctrl.c2d_rf_waddr_W[0] ),
    .B1(_02091_),
    .C1(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__or4b_4 _07878_ (.A(_02086_),
    .B(_02090_),
    .C(_02093_),
    .D_N(_01981_),
    .X(_02094_));
 sky130_fd_sc_hd__and2_4 _07879_ (.A(_02001_),
    .B(_02076_),
    .X(_02095_));
 sky130_fd_sc_hd__a21bo_1 _07880_ (.A1(_02001_),
    .A2(_02076_),
    .B1_N(_02062_),
    .X(_02096_));
 sky130_fd_sc_hd__nand2b_4 _07881_ (.A_N(_02096_),
    .B(_02094_),
    .Y(_02097_));
 sky130_fd_sc_hd__nor3_1 _07882_ (.A(_02052_),
    .B(net482),
    .C(net372),
    .Y(_02098_));
 sky130_fd_sc_hd__mux2_4 _07883_ (.A0(net3589),
    .A1(net23),
    .S(net480),
    .X(_02099_));
 sky130_fd_sc_hd__and2_2 _07884_ (.A(_01961_),
    .B(_02067_),
    .X(_02100_));
 sky130_fd_sc_hd__nand2_4 _07885_ (.A(_01961_),
    .B(_02067_),
    .Y(_02101_));
 sky130_fd_sc_hd__a21oi_1 _07886_ (.A1(_01842_),
    .A2(_01905_),
    .B1(_01904_),
    .Y(_02102_));
 sky130_fd_sc_hd__xnor2_1 _07887_ (.A(_01857_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__a21o_1 _07888_ (.A1(net651),
    .A2(net780),
    .B1(_01904_),
    .X(_02104_));
 sky130_fd_sc_hd__nand3_2 _07889_ (.A(net651),
    .B(net780),
    .C(_01904_),
    .Y(_02105_));
 sky130_fd_sc_hd__nand4_2 _07890_ (.A(net786),
    .B(net643),
    .C(_02104_),
    .D(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__a22o_1 _07891_ (.A1(net786),
    .A2(net643),
    .B1(_02104_),
    .B2(_02105_),
    .X(_02107_));
 sky130_fd_sc_hd__and4_1 _07892_ (.A(net651),
    .B(net786),
    .C(net647),
    .D(net783),
    .X(_02108_));
 sky130_fd_sc_hd__a21oi_1 _07893_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__and3_1 _07894_ (.A(_02106_),
    .B(_02107_),
    .C(_02108_),
    .X(_02110_));
 sky130_fd_sc_hd__inv_2 _07895_ (.A(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__o21ai_1 _07896_ (.A1(_02109_),
    .A2(_02110_),
    .B1(net484),
    .Y(_02112_));
 sky130_fd_sc_hd__o211a_1 _07897_ (.A1(net3684),
    .A2(net484),
    .B1(net468),
    .C1(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__a21o_4 _07898_ (.A1(net467),
    .A2(_02103_),
    .B1(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__nor2_2 _07899_ (.A(_02094_),
    .B(_02096_),
    .Y(_02115_));
 sky130_fd_sc_hd__nor2_2 _07900_ (.A(_02062_),
    .B(net392),
    .Y(_02116_));
 sky130_fd_sc_hd__a22o_1 _07901_ (.A1(net392),
    .A2(_02114_),
    .B1(net368),
    .B2(_02099_),
    .X(_02117_));
 sky130_fd_sc_hd__a211o_2 _07902_ (.A1(net714),
    .A2(net370),
    .B1(_02117_),
    .C1(_02098_),
    .X(_02118_));
 sky130_fd_sc_hd__nand3b_2 _07903_ (.A_N(net404),
    .B(_01836_),
    .C(net3465),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_2 _07904_ (.A(_01974_),
    .B(_01982_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21o_1 _07905_ (.A1(_01974_),
    .A2(_01982_),
    .B1(net3235),
    .X(_02121_));
 sky130_fd_sc_hd__or3b_1 _07906_ (.A(net3393),
    .B(_01973_),
    .C_N(_01982_),
    .X(_02122_));
 sky130_fd_sc_hd__and2_1 _07907_ (.A(_02121_),
    .B(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__and3_1 _07908_ (.A(net3233),
    .B(_02121_),
    .C(_02122_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_2 _07909_ (.A(_01836_),
    .B(_01973_),
    .Y(_02125_));
 sky130_fd_sc_hd__or2_2 _07910_ (.A(_01836_),
    .B(_01973_),
    .X(_02126_));
 sky130_fd_sc_hd__a21o_1 _07911_ (.A1(_01974_),
    .A2(_01982_),
    .B1(net3205),
    .X(_02127_));
 sky130_fd_sc_hd__o21a_1 _07912_ (.A1(net3432),
    .A2(_02120_),
    .B1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__o2111a_1 _07913_ (.A1(net3432),
    .A2(_02120_),
    .B1(_02125_),
    .C1(_02127_),
    .D1(net3249),
    .X(_02129_));
 sky130_fd_sc_hd__a21o_1 _07914_ (.A1(_02121_),
    .A2(_02122_),
    .B1(net3233),
    .X(_02130_));
 sky130_fd_sc_hd__nand2b_1 _07915_ (.A_N(_02124_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21o_1 _07916_ (.A1(_02129_),
    .A2(_02130_),
    .B1(_02124_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_2 _07917_ (.A0(net3403),
    .A1(net3202),
    .S(_02120_),
    .X(_02133_));
 sky130_fd_sc_hd__or2_1 _07918_ (.A(net3518),
    .B(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(net3518),
    .B(_02133_),
    .Y(_02135_));
 sky130_fd_sc_hd__and2_1 _07920_ (.A(_02134_),
    .B(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__xnor2_1 _07921_ (.A(_02132_),
    .B(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _07922_ (.A(net366),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_1 _07923_ (.A(net250),
    .B(net443),
    .Y(_02139_));
 sky130_fd_sc_hd__a211o_1 _07924_ (.A1(net250),
    .A2(net444),
    .B1(_02010_),
    .C1(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__a221o_1 _07925_ (.A1(net3475),
    .A2(net404),
    .B1(_02027_),
    .B2(_02118_),
    .C1(_02138_),
    .X(_02141_));
 sky130_fd_sc_hd__nand2_1 _07926_ (.A(_02010_),
    .B(net3476),
    .Y(_02142_));
 sky130_fd_sc_hd__a21oi_1 _07927_ (.A1(_02140_),
    .A2(_02142_),
    .B1(net880),
    .Y(_00638_));
 sky130_fd_sc_hd__mux4_1 _07928_ (.A0(\dpath.RF.R[0][3] ),
    .A1(\dpath.RF.R[1][3] ),
    .A2(\dpath.RF.R[2][3] ),
    .A3(\dpath.RF.R[3][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02143_));
 sky130_fd_sc_hd__mux4_1 _07929_ (.A0(\dpath.RF.R[4][3] ),
    .A1(\dpath.RF.R[5][3] ),
    .A2(\dpath.RF.R[6][3] ),
    .A3(\dpath.RF.R[7][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02144_));
 sky130_fd_sc_hd__o21a_1 _07930_ (.A1(net508),
    .A2(_02144_),
    .B1(net506),
    .X(_02145_));
 sky130_fd_sc_hd__o21ai_1 _07931_ (.A1(net529),
    .A2(_02143_),
    .B1(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__mux4_1 _07932_ (.A0(\dpath.RF.R[12][3] ),
    .A1(\dpath.RF.R[13][3] ),
    .A2(\dpath.RF.R[14][3] ),
    .A3(\dpath.RF.R[15][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02147_));
 sky130_fd_sc_hd__mux4_1 _07933_ (.A0(\dpath.RF.R[8][3] ),
    .A1(\dpath.RF.R[9][3] ),
    .A2(\dpath.RF.R[10][3] ),
    .A3(\dpath.RF.R[11][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02148_));
 sky130_fd_sc_hd__or2_1 _07934_ (.A(net529),
    .B(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__o211a_1 _07935_ (.A1(net508),
    .A2(_02147_),
    .B1(_02149_),
    .C1(net521),
    .X(_02150_));
 sky130_fd_sc_hd__nor2_1 _07936_ (.A(net517),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__mux4_1 _07937_ (.A0(\dpath.RF.R[16][3] ),
    .A1(\dpath.RF.R[17][3] ),
    .A2(\dpath.RF.R[18][3] ),
    .A3(\dpath.RF.R[19][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02152_));
 sky130_fd_sc_hd__nor2_1 _07938_ (.A(net529),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__mux4_1 _07939_ (.A0(\dpath.RF.R[20][3] ),
    .A1(\dpath.RF.R[21][3] ),
    .A2(\dpath.RF.R[22][3] ),
    .A3(\dpath.RF.R[23][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02154_));
 sky130_fd_sc_hd__nor2_1 _07940_ (.A(net508),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__mux4_1 _07941_ (.A0(\dpath.RF.R[28][3] ),
    .A1(\dpath.RF.R[29][3] ),
    .A2(\dpath.RF.R[30][3] ),
    .A3(\dpath.RF.R[31][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02156_));
 sky130_fd_sc_hd__nor2_1 _07942_ (.A(net508),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__mux4_1 _07943_ (.A0(\dpath.RF.R[24][3] ),
    .A1(\dpath.RF.R[25][3] ),
    .A2(\dpath.RF.R[26][3] ),
    .A3(\dpath.RF.R[27][3] ),
    .S0(net557),
    .S1(net538),
    .X(_02158_));
 sky130_fd_sc_hd__o21ai_1 _07944_ (.A1(net529),
    .A2(_02158_),
    .B1(net521),
    .Y(_02159_));
 sky130_fd_sc_hd__o32a_1 _07945_ (.A1(net521),
    .A2(_02153_),
    .A3(_02155_),
    .B1(_02157_),
    .B2(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__a221o_1 _07946_ (.A1(_02146_),
    .A2(_02151_),
    .B1(_02160_),
    .B2(net517),
    .C1(net482),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_1 _07947_ (.A(net372),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__mux2_1 _07948_ (.A0(net3650),
    .A1(net26),
    .S(net480),
    .X(_02163_));
 sky130_fd_sc_hd__a221o_1 _07949_ (.A1(net713),
    .A2(net370),
    .B1(net368),
    .B2(_02163_),
    .C1(_02162_),
    .X(_02164_));
 sky130_fd_sc_hd__o21ai_1 _07950_ (.A1(_01856_),
    .A2(_02102_),
    .B1(_01854_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_1 _07951_ (.A(_01903_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__a22oi_1 _07952_ (.A1(net647),
    .A2(net780),
    .B1(net776),
    .B2(net651),
    .Y(_02167_));
 sky130_fd_sc_hd__and4_1 _07953_ (.A(net651),
    .B(net647),
    .C(net780),
    .D(net776),
    .X(_02168_));
 sky130_fd_sc_hd__and4bb_1 _07954_ (.A_N(_02167_),
    .B_N(_02168_),
    .C(net783),
    .D(net643),
    .X(_02169_));
 sky130_fd_sc_hd__o2bb2a_1 _07955_ (.A1_N(net783),
    .A2_N(net643),
    .B1(_02167_),
    .B2(_02168_),
    .X(_02170_));
 sky130_fd_sc_hd__or2_1 _07956_ (.A(_02169_),
    .B(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__or2_1 _07957_ (.A(_02105_),
    .B(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__nand2_1 _07958_ (.A(_02105_),
    .B(_02171_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(_02172_),
    .B(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand2_1 _07960_ (.A(net786),
    .B(net638),
    .Y(_02175_));
 sky130_fd_sc_hd__xnor2_1 _07961_ (.A(_02174_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _07962_ (.A(_02106_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__and2_1 _07963_ (.A(_02106_),
    .B(_02176_),
    .X(_02178_));
 sky130_fd_sc_hd__or2_1 _07964_ (.A(_02177_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__nor2_1 _07965_ (.A(_02111_),
    .B(_02176_),
    .Y(_02180_));
 sky130_fd_sc_hd__a21oi_1 _07966_ (.A1(_02111_),
    .A2(_02179_),
    .B1(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__mux2_1 _07967_ (.A0(net3683),
    .A1(_02181_),
    .S(net484),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_4 _07968_ (.A0(_02166_),
    .A1(_02182_),
    .S(net468),
    .X(_02183_));
 sky130_fd_sc_hd__a21oi_1 _07969_ (.A1(net392),
    .A2(_02183_),
    .B1(net3272),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _07970_ (.A(net373),
    .B(net3273),
    .Y(_02185_));
 sky130_fd_sc_hd__a21bo_1 _07971_ (.A1(_02132_),
    .A2(_02134_),
    .B1_N(_02135_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_2 _07972_ (.A0(net3285),
    .A1(net3237),
    .S(_02120_),
    .X(_02187_));
 sky130_fd_sc_hd__or2_1 _07973_ (.A(net3231),
    .B(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(net3231),
    .B(_02187_),
    .Y(_02189_));
 sky130_fd_sc_hd__and2_1 _07975_ (.A(_02188_),
    .B(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__xnor2_1 _07976_ (.A(_02186_),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _07977_ (.A(net366),
    .B(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_1 _07978_ (.A(net3493),
    .B(net250),
    .Y(_02193_));
 sky130_fd_sc_hd__or2_1 _07979_ (.A(net3493),
    .B(net250),
    .X(_02194_));
 sky130_fd_sc_hd__a32o_1 _07980_ (.A1(net362),
    .A2(_02193_),
    .A3(_02194_),
    .B1(net403),
    .B2(\dpath.btarg_DX.q[3] ),
    .X(_02195_));
 sky130_fd_sc_hd__or3_1 _07981_ (.A(_02008_),
    .B(_02192_),
    .C(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__o221a_1 _07982_ (.A1(net3493),
    .A2(net444),
    .B1(_02185_),
    .B2(_02196_),
    .C1(net843),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_1 _07983_ (.A0(\dpath.RF.R[0][4] ),
    .A1(\dpath.RF.R[1][4] ),
    .A2(\dpath.RF.R[2][4] ),
    .A3(\dpath.RF.R[3][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02197_));
 sky130_fd_sc_hd__mux4_1 _07984_ (.A0(\dpath.RF.R[4][4] ),
    .A1(\dpath.RF.R[5][4] ),
    .A2(\dpath.RF.R[6][4] ),
    .A3(\dpath.RF.R[7][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02198_));
 sky130_fd_sc_hd__o21a_1 _07985_ (.A1(net508),
    .A2(_02198_),
    .B1(net506),
    .X(_02199_));
 sky130_fd_sc_hd__o21ai_1 _07986_ (.A1(net529),
    .A2(_02197_),
    .B1(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__mux4_1 _07987_ (.A0(\dpath.RF.R[12][4] ),
    .A1(\dpath.RF.R[13][4] ),
    .A2(\dpath.RF.R[14][4] ),
    .A3(\dpath.RF.R[15][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02201_));
 sky130_fd_sc_hd__mux4_1 _07988_ (.A0(\dpath.RF.R[8][4] ),
    .A1(\dpath.RF.R[9][4] ),
    .A2(\dpath.RF.R[10][4] ),
    .A3(\dpath.RF.R[11][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02202_));
 sky130_fd_sc_hd__or2_1 _07989_ (.A(net529),
    .B(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__o211a_1 _07990_ (.A1(net508),
    .A2(_02201_),
    .B1(_02203_),
    .C1(net521),
    .X(_02204_));
 sky130_fd_sc_hd__nor2_1 _07991_ (.A(net517),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__mux4_1 _07992_ (.A0(\dpath.RF.R[16][4] ),
    .A1(\dpath.RF.R[17][4] ),
    .A2(\dpath.RF.R[18][4] ),
    .A3(\dpath.RF.R[19][4] ),
    .S0(net561),
    .S1(net542),
    .X(_02206_));
 sky130_fd_sc_hd__nor2_1 _07993_ (.A(net529),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__mux4_1 _07994_ (.A0(\dpath.RF.R[20][4] ),
    .A1(\dpath.RF.R[21][4] ),
    .A2(\dpath.RF.R[22][4] ),
    .A3(\dpath.RF.R[23][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02208_));
 sky130_fd_sc_hd__nor2_1 _07995_ (.A(net510),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__mux4_1 _07996_ (.A0(\dpath.RF.R[28][4] ),
    .A1(\dpath.RF.R[29][4] ),
    .A2(\dpath.RF.R[30][4] ),
    .A3(\dpath.RF.R[31][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02210_));
 sky130_fd_sc_hd__nor2_1 _07997_ (.A(net510),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__mux4_1 _07998_ (.A0(\dpath.RF.R[24][4] ),
    .A1(\dpath.RF.R[25][4] ),
    .A2(\dpath.RF.R[26][4] ),
    .A3(\dpath.RF.R[27][4] ),
    .S0(net558),
    .S1(net539),
    .X(_02212_));
 sky130_fd_sc_hd__o21ai_1 _07999_ (.A1(net529),
    .A2(_02212_),
    .B1(net521),
    .Y(_02213_));
 sky130_fd_sc_hd__o32a_1 _08000_ (.A1(net521),
    .A2(_02207_),
    .A3(_02209_),
    .B1(_02211_),
    .B2(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__a221o_1 _08001_ (.A1(_02200_),
    .A2(_02205_),
    .B1(_02214_),
    .B2(net517),
    .C1(net482),
    .X(_02215_));
 sky130_fd_sc_hd__nor2_1 _08002_ (.A(net372),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__mux2_2 _08003_ (.A0(net3651),
    .A1(net27),
    .S(net480),
    .X(_02217_));
 sky130_fd_sc_hd__a221o_1 _08004_ (.A1(net3267),
    .A2(net370),
    .B1(net368),
    .B2(_02217_),
    .C1(_02216_),
    .X(_02218_));
 sky130_fd_sc_hd__and4_1 _08005_ (.A(net651),
    .B(net647),
    .C(net776),
    .D(net772),
    .X(_02219_));
 sky130_fd_sc_hd__a22oi_2 _08006_ (.A1(net647),
    .A2(net776),
    .B1(net772),
    .B2(net651),
    .Y(_02220_));
 sky130_fd_sc_hd__or3_1 _08007_ (.A(_01854_),
    .B(_02219_),
    .C(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__o21ai_1 _08008_ (.A1(_02219_),
    .A2(_02220_),
    .B1(_01854_),
    .Y(_02222_));
 sky130_fd_sc_hd__and3_1 _08009_ (.A(_02168_),
    .B(_02221_),
    .C(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__nand3_1 _08010_ (.A(_02168_),
    .B(_02221_),
    .C(_02222_),
    .Y(_02224_));
 sky130_fd_sc_hd__a21o_1 _08011_ (.A1(_02221_),
    .A2(_02222_),
    .B1(_02168_),
    .X(_02225_));
 sky130_fd_sc_hd__nand4_1 _08012_ (.A(net783),
    .B(net638),
    .C(_02224_),
    .D(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__a22o_1 _08013_ (.A1(net783),
    .A2(net638),
    .B1(_02224_),
    .B2(_02225_),
    .X(_02227_));
 sky130_fd_sc_hd__nand3_1 _08014_ (.A(_02169_),
    .B(_02226_),
    .C(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__a21o_1 _08015_ (.A1(_02226_),
    .A2(_02227_),
    .B1(_02169_),
    .X(_02229_));
 sky130_fd_sc_hd__and2_1 _08016_ (.A(net786),
    .B(\dpath.alu.adder.in0[4] ),
    .X(_02230_));
 sky130_fd_sc_hd__nand3_1 _08017_ (.A(_02228_),
    .B(_02229_),
    .C(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__a21o_1 _08018_ (.A1(_02228_),
    .A2(_02229_),
    .B1(_02230_),
    .X(_02232_));
 sky130_fd_sc_hd__o21ai_1 _08019_ (.A1(_02174_),
    .A2(_02175_),
    .B1(_02172_),
    .Y(_02233_));
 sky130_fd_sc_hd__and3_1 _08020_ (.A(_02231_),
    .B(_02232_),
    .C(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__a21oi_1 _08021_ (.A1(_02231_),
    .A2(_02232_),
    .B1(_02233_),
    .Y(_02235_));
 sky130_fd_sc_hd__nor3b_1 _08022_ (.A(_02234_),
    .B(_02235_),
    .C_N(_02177_),
    .Y(_02236_));
 sky130_fd_sc_hd__o21bai_1 _08023_ (.A1(_02234_),
    .A2(_02235_),
    .B1_N(_02177_),
    .Y(_02237_));
 sky130_fd_sc_hd__and2b_1 _08024_ (.A_N(_02236_),
    .B(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__nor2_4 _08025_ (.A(net485),
    .B(net467),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_8 _08026_ (.A(net484),
    .B(net468),
    .Y(_02240_));
 sky130_fd_sc_hd__a21oi_1 _08027_ (.A1(_02180_),
    .A2(_02238_),
    .B1(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__o21a_1 _08028_ (.A1(_02180_),
    .A2(_02238_),
    .B1(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__a21bo_1 _08029_ (.A1(_01901_),
    .A2(_02165_),
    .B1_N(_01902_),
    .X(_02243_));
 sky130_fd_sc_hd__a21oi_1 _08030_ (.A1(_01853_),
    .A2(_02243_),
    .B1(net468),
    .Y(_02244_));
 sky130_fd_sc_hd__o21a_1 _08031_ (.A1(_01853_),
    .A2(_02243_),
    .B1(_02244_),
    .X(_02245_));
 sky130_fd_sc_hd__a211o_4 _08032_ (.A1(net3543),
    .A2(net485),
    .B1(_02242_),
    .C1(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__a21oi_1 _08033_ (.A1(net392),
    .A2(_02246_),
    .B1(net3268),
    .Y(_02247_));
 sky130_fd_sc_hd__nor2_1 _08034_ (.A(net373),
    .B(net3269),
    .Y(_02248_));
 sky130_fd_sc_hd__a21bo_1 _08035_ (.A1(_02186_),
    .A2(_02188_),
    .B1_N(_02189_),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_2 _08036_ (.A0(net3349),
    .A1(net3219),
    .S(_02120_),
    .X(_02250_));
 sky130_fd_sc_hd__or2_1 _08037_ (.A(net3238),
    .B(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__nand2_1 _08038_ (.A(net3238),
    .B(_02250_),
    .Y(_02252_));
 sky130_fd_sc_hd__and2_1 _08039_ (.A(_02251_),
    .B(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__xnor2_1 _08040_ (.A(_02249_),
    .B(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _08041_ (.A(net365),
    .B(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__and3_1 _08042_ (.A(net254),
    .B(net3493),
    .C(net250),
    .X(_02256_));
 sky130_fd_sc_hd__inv_2 _08043_ (.A(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__a21o_1 _08044_ (.A1(net253),
    .A2(net250),
    .B1(net254),
    .X(_02258_));
 sky130_fd_sc_hd__a32o_1 _08045_ (.A1(net361),
    .A2(_02257_),
    .A3(_02258_),
    .B1(net403),
    .B2(net3478),
    .X(_02259_));
 sky130_fd_sc_hd__or3_1 _08046_ (.A(net450),
    .B(_02255_),
    .C(net3479),
    .X(_02260_));
 sky130_fd_sc_hd__o221a_1 _08047_ (.A1(net254),
    .A2(net442),
    .B1(_02248_),
    .B2(_02260_),
    .C1(net846),
    .X(_00640_));
 sky130_fd_sc_hd__and2_1 _08048_ (.A(net3280),
    .B(_02256_),
    .X(_02261_));
 sky130_fd_sc_hd__nor2_1 _08049_ (.A(net3280),
    .B(_02256_),
    .Y(_02262_));
 sky130_fd_sc_hd__o21a_1 _08050_ (.A1(_02261_),
    .A2(_02262_),
    .B1(net361),
    .X(_02263_));
 sky130_fd_sc_hd__mux4_1 _08051_ (.A0(\dpath.RF.R[0][5] ),
    .A1(\dpath.RF.R[1][5] ),
    .A2(\dpath.RF.R[2][5] ),
    .A3(\dpath.RF.R[3][5] ),
    .S0(net558),
    .S1(net539),
    .X(_02264_));
 sky130_fd_sc_hd__mux4_1 _08052_ (.A0(\dpath.RF.R[4][5] ),
    .A1(\dpath.RF.R[5][5] ),
    .A2(\dpath.RF.R[6][5] ),
    .A3(\dpath.RF.R[7][5] ),
    .S0(net558),
    .S1(net539),
    .X(_02265_));
 sky130_fd_sc_hd__o21a_1 _08053_ (.A1(net508),
    .A2(_02265_),
    .B1(net506),
    .X(_02266_));
 sky130_fd_sc_hd__o21ai_1 _08054_ (.A1(net529),
    .A2(_02264_),
    .B1(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__mux4_1 _08055_ (.A0(\dpath.RF.R[12][5] ),
    .A1(\dpath.RF.R[13][5] ),
    .A2(\dpath.RF.R[14][5] ),
    .A3(\dpath.RF.R[15][5] ),
    .S0(net560),
    .S1(net541),
    .X(_02268_));
 sky130_fd_sc_hd__mux4_1 _08056_ (.A0(\dpath.RF.R[8][5] ),
    .A1(\dpath.RF.R[9][5] ),
    .A2(\dpath.RF.R[10][5] ),
    .A3(\dpath.RF.R[11][5] ),
    .S0(net560),
    .S1(net541),
    .X(_02269_));
 sky130_fd_sc_hd__or2_1 _08057_ (.A(net530),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__o211a_1 _08058_ (.A1(net510),
    .A2(_02268_),
    .B1(_02270_),
    .C1(net522),
    .X(_02271_));
 sky130_fd_sc_hd__nor2_1 _08059_ (.A(net517),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__mux4_1 _08060_ (.A0(\dpath.RF.R[16][5] ),
    .A1(\dpath.RF.R[17][5] ),
    .A2(\dpath.RF.R[18][5] ),
    .A3(\dpath.RF.R[19][5] ),
    .S0(net560),
    .S1(net541),
    .X(_02273_));
 sky130_fd_sc_hd__nor2_1 _08061_ (.A(net530),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__mux4_1 _08062_ (.A0(\dpath.RF.R[20][5] ),
    .A1(\dpath.RF.R[21][5] ),
    .A2(\dpath.RF.R[22][5] ),
    .A3(\dpath.RF.R[23][5] ),
    .S0(net558),
    .S1(net539),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_1 _08063_ (.A(net508),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__mux4_1 _08064_ (.A0(\dpath.RF.R[28][5] ),
    .A1(\dpath.RF.R[29][5] ),
    .A2(\dpath.RF.R[30][5] ),
    .A3(\dpath.RF.R[31][5] ),
    .S0(net560),
    .S1(net541),
    .X(_02277_));
 sky130_fd_sc_hd__nor2_1 _08065_ (.A(net510),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__mux4_1 _08066_ (.A0(\dpath.RF.R[24][5] ),
    .A1(\dpath.RF.R[25][5] ),
    .A2(\dpath.RF.R[26][5] ),
    .A3(\dpath.RF.R[27][5] ),
    .S0(net560),
    .S1(net541),
    .X(_02279_));
 sky130_fd_sc_hd__o21ai_1 _08067_ (.A1(net533),
    .A2(_02279_),
    .B1(net521),
    .Y(_02280_));
 sky130_fd_sc_hd__o32a_1 _08068_ (.A1(net521),
    .A2(_02274_),
    .A3(_02276_),
    .B1(_02278_),
    .B2(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__a221o_1 _08069_ (.A1(_02267_),
    .A2(_02272_),
    .B1(_02281_),
    .B2(net517),
    .C1(net482),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_1 _08070_ (.A(net372),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__mux2_2 _08071_ (.A0(net3624),
    .A1(net28),
    .S(net480),
    .X(_02284_));
 sky130_fd_sc_hd__a221o_1 _08072_ (.A1(net708),
    .A2(net370),
    .B1(net368),
    .B2(_02284_),
    .C1(_02283_),
    .X(_02285_));
 sky130_fd_sc_hd__nand2_1 _08073_ (.A(net783),
    .B(net632),
    .Y(_02286_));
 sky130_fd_sc_hd__and2_1 _08074_ (.A(net780),
    .B(net636),
    .X(_02287_));
 sky130_fd_sc_hd__nand4_2 _08075_ (.A(net647),
    .B(net643),
    .C(net776),
    .D(net772),
    .Y(_02288_));
 sky130_fd_sc_hd__a22o_1 _08076_ (.A1(net643),
    .A2(net776),
    .B1(net772),
    .B2(net647),
    .X(_02289_));
 sky130_fd_sc_hd__nand3_1 _08077_ (.A(_02287_),
    .B(_02288_),
    .C(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__a21o_1 _08078_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02287_),
    .X(_02291_));
 sky130_fd_sc_hd__o21bai_1 _08079_ (.A1(_01854_),
    .A2(_02220_),
    .B1_N(_02219_),
    .Y(_02292_));
 sky130_fd_sc_hd__and3_1 _08080_ (.A(_02290_),
    .B(_02291_),
    .C(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__a21oi_1 _08081_ (.A1(_02290_),
    .A2(_02291_),
    .B1(_02292_),
    .Y(_02294_));
 sky130_fd_sc_hd__or3_1 _08082_ (.A(_02286_),
    .B(_02293_),
    .C(_02294_),
    .X(_02295_));
 sky130_fd_sc_hd__o21ai_1 _08083_ (.A1(_02293_),
    .A2(_02294_),
    .B1(_02286_),
    .Y(_02296_));
 sky130_fd_sc_hd__a31o_1 _08084_ (.A1(net783),
    .A2(net638),
    .A3(_02225_),
    .B1(_02223_),
    .X(_02297_));
 sky130_fd_sc_hd__nand3_1 _08085_ (.A(_02295_),
    .B(_02296_),
    .C(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__a21o_1 _08086_ (.A1(_02295_),
    .A2(_02296_),
    .B1(_02297_),
    .X(_02299_));
 sky130_fd_sc_hd__a22o_1 _08087_ (.A1(net786),
    .A2(net628),
    .B1(_02298_),
    .B2(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__nand4_2 _08088_ (.A(net786),
    .B(net628),
    .C(_02298_),
    .D(_02299_),
    .Y(_02301_));
 sky130_fd_sc_hd__and4_2 _08089_ (.A(net651),
    .B(net768),
    .C(_02300_),
    .D(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__a22oi_2 _08090_ (.A1(net651),
    .A2(net768),
    .B1(_02300_),
    .B2(_02301_),
    .Y(_02303_));
 sky130_fd_sc_hd__and2_1 _08091_ (.A(_02228_),
    .B(_02231_),
    .X(_02304_));
 sky130_fd_sc_hd__nor3_1 _08092_ (.A(_02302_),
    .B(_02303_),
    .C(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__or3_1 _08093_ (.A(_02302_),
    .B(_02303_),
    .C(_02304_),
    .X(_02306_));
 sky130_fd_sc_hd__o21ai_1 _08094_ (.A1(_02302_),
    .A2(_02303_),
    .B1(_02304_),
    .Y(_02307_));
 sky130_fd_sc_hd__and3_1 _08095_ (.A(_02234_),
    .B(_02306_),
    .C(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__a21oi_1 _08096_ (.A1(_02306_),
    .A2(_02307_),
    .B1(_02234_),
    .Y(_02309_));
 sky130_fd_sc_hd__or2_1 _08097_ (.A(_02308_),
    .B(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__a21oi_2 _08098_ (.A1(_02180_),
    .A2(_02237_),
    .B1(_02236_),
    .Y(_02311_));
 sky130_fd_sc_hd__a21oi_1 _08099_ (.A1(_02310_),
    .A2(_02311_),
    .B1(_02240_),
    .Y(_02312_));
 sky130_fd_sc_hd__o21a_1 _08100_ (.A1(_02310_),
    .A2(_02311_),
    .B1(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__a21oi_1 _08101_ (.A1(_01853_),
    .A2(_02243_),
    .B1(_01851_),
    .Y(_02314_));
 sky130_fd_sc_hd__xnor2_1 _08102_ (.A(_01847_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__a221o_4 _08103_ (.A1(net3653),
    .A2(net485),
    .B1(net467),
    .B2(_02315_),
    .C1(_02313_),
    .X(_02316_));
 sky130_fd_sc_hd__a21oi_4 _08104_ (.A1(net392),
    .A2(_02316_),
    .B1(_02285_),
    .Y(_02317_));
 sky130_fd_sc_hd__a21boi_1 _08105_ (.A1(_02249_),
    .A2(_02251_),
    .B1_N(_02252_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_1 _08106_ (.A(net3392),
    .B(net1338),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _08107_ (.A(net3392),
    .B(net1338),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2b_1 _08108_ (.A_N(_02319_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_1 _08109_ (.A(_02318_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__a21oi_1 _08110_ (.A1(net3534),
    .A2(net403),
    .B1(net361),
    .Y(_02323_));
 sky130_fd_sc_hd__o221a_1 _08111_ (.A1(net373),
    .A2(_02317_),
    .B1(_02322_),
    .B2(net365),
    .C1(_02323_),
    .X(_02324_));
 sky130_fd_sc_hd__o21ai_1 _08112_ (.A1(_02263_),
    .A2(_02324_),
    .B1(net442),
    .Y(_02325_));
 sky130_fd_sc_hd__o211a_1 _08113_ (.A1(net3280),
    .A2(net442),
    .B1(net3535),
    .C1(net846),
    .X(_00641_));
 sky130_fd_sc_hd__xnor2_1 _08114_ (.A(net256),
    .B(_02261_),
    .Y(_02326_));
 sky130_fd_sc_hd__mux4_1 _08115_ (.A0(\dpath.RF.R[0][6] ),
    .A1(\dpath.RF.R[1][6] ),
    .A2(\dpath.RF.R[2][6] ),
    .A3(\dpath.RF.R[3][6] ),
    .S0(net558),
    .S1(net539),
    .X(_02327_));
 sky130_fd_sc_hd__mux4_1 _08116_ (.A0(\dpath.RF.R[4][6] ),
    .A1(\dpath.RF.R[5][6] ),
    .A2(\dpath.RF.R[6][6] ),
    .A3(\dpath.RF.R[7][6] ),
    .S0(net558),
    .S1(net539),
    .X(_02328_));
 sky130_fd_sc_hd__o21a_1 _08117_ (.A1(net510),
    .A2(_02328_),
    .B1(net506),
    .X(_02329_));
 sky130_fd_sc_hd__o21ai_1 _08118_ (.A1(net533),
    .A2(_02327_),
    .B1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__mux4_1 _08119_ (.A0(\dpath.RF.R[12][6] ),
    .A1(\dpath.RF.R[13][6] ),
    .A2(\dpath.RF.R[14][6] ),
    .A3(\dpath.RF.R[15][6] ),
    .S0(net558),
    .S1(net539),
    .X(_02331_));
 sky130_fd_sc_hd__mux4_1 _08120_ (.A0(\dpath.RF.R[8][6] ),
    .A1(\dpath.RF.R[9][6] ),
    .A2(\dpath.RF.R[10][6] ),
    .A3(\dpath.RF.R[11][6] ),
    .S0(net558),
    .S1(net539),
    .X(_02332_));
 sky130_fd_sc_hd__or2_1 _08121_ (.A(net529),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__o211a_1 _08122_ (.A1(net508),
    .A2(_02331_),
    .B1(_02333_),
    .C1(net521),
    .X(_02334_));
 sky130_fd_sc_hd__nor2_1 _08123_ (.A(net517),
    .B(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__mux4_1 _08124_ (.A0(\dpath.RF.R[16][6] ),
    .A1(\dpath.RF.R[17][6] ),
    .A2(\dpath.RF.R[18][6] ),
    .A3(\dpath.RF.R[19][6] ),
    .S0(net562),
    .S1(net543),
    .X(_02336_));
 sky130_fd_sc_hd__nor2_1 _08125_ (.A(net533),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__mux4_1 _08126_ (.A0(\dpath.RF.R[20][6] ),
    .A1(\dpath.RF.R[21][6] ),
    .A2(\dpath.RF.R[22][6] ),
    .A3(\dpath.RF.R[23][6] ),
    .S0(net558),
    .S1(net539),
    .X(_02338_));
 sky130_fd_sc_hd__nor2_1 _08127_ (.A(net508),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__mux4_1 _08128_ (.A0(\dpath.RF.R[28][6] ),
    .A1(\dpath.RF.R[29][6] ),
    .A2(\dpath.RF.R[30][6] ),
    .A3(\dpath.RF.R[31][6] ),
    .S0(net561),
    .S1(net542),
    .X(_02340_));
 sky130_fd_sc_hd__nor2_1 _08129_ (.A(net508),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__mux4_1 _08130_ (.A0(\dpath.RF.R[24][6] ),
    .A1(\dpath.RF.R[25][6] ),
    .A2(\dpath.RF.R[26][6] ),
    .A3(\dpath.RF.R[27][6] ),
    .S0(net558),
    .S1(net539),
    .X(_02342_));
 sky130_fd_sc_hd__o21ai_1 _08131_ (.A1(net529),
    .A2(_02342_),
    .B1(net521),
    .Y(_02343_));
 sky130_fd_sc_hd__o32a_1 _08132_ (.A1(net521),
    .A2(_02337_),
    .A3(_02339_),
    .B1(_02341_),
    .B2(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__a221o_1 _08133_ (.A1(_02330_),
    .A2(_02335_),
    .B1(_02344_),
    .B2(net517),
    .C1(net482),
    .X(_02345_));
 sky130_fd_sc_hd__nor2_1 _08134_ (.A(net372),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__mux2_2 _08135_ (.A0(net3411),
    .A1(net29),
    .S(net480),
    .X(_02347_));
 sky130_fd_sc_hd__a221o_1 _08136_ (.A1(net707),
    .A2(net370),
    .B1(net368),
    .B2(_02347_),
    .C1(_02346_),
    .X(_02348_));
 sky130_fd_sc_hd__a22oi_1 _08137_ (.A1(net646),
    .A2(net770),
    .B1(net765),
    .B2(net650),
    .Y(_02349_));
 sky130_fd_sc_hd__and4_1 _08138_ (.A(net650),
    .B(net646),
    .C(net770),
    .D(net765),
    .X(_02350_));
 sky130_fd_sc_hd__nor2_1 _08139_ (.A(_02349_),
    .B(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2_1 _08140_ (.A(net783),
    .B(net628),
    .Y(_02352_));
 sky130_fd_sc_hd__and2_1 _08141_ (.A(net780),
    .B(net632),
    .X(_02353_));
 sky130_fd_sc_hd__nand4_1 _08142_ (.A(net641),
    .B(net636),
    .C(net776),
    .D(net772),
    .Y(_02354_));
 sky130_fd_sc_hd__a22o_1 _08143_ (.A1(net636),
    .A2(net776),
    .B1(net772),
    .B2(net641),
    .X(_02355_));
 sky130_fd_sc_hd__nand3_1 _08144_ (.A(_02353_),
    .B(_02354_),
    .C(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__a21o_1 _08145_ (.A1(_02354_),
    .A2(_02355_),
    .B1(_02353_),
    .X(_02357_));
 sky130_fd_sc_hd__a21bo_1 _08146_ (.A1(_02287_),
    .A2(_02289_),
    .B1_N(_02288_),
    .X(_02358_));
 sky130_fd_sc_hd__and3_1 _08147_ (.A(_02356_),
    .B(_02357_),
    .C(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__a21oi_1 _08148_ (.A1(_02356_),
    .A2(_02357_),
    .B1(_02358_),
    .Y(_02360_));
 sky130_fd_sc_hd__or3_1 _08149_ (.A(_02352_),
    .B(_02359_),
    .C(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__o21ai_1 _08150_ (.A1(_02359_),
    .A2(_02360_),
    .B1(_02352_),
    .Y(_02362_));
 sky130_fd_sc_hd__o21bai_2 _08151_ (.A1(_02286_),
    .A2(_02294_),
    .B1_N(_02293_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand3_2 _08152_ (.A(_02361_),
    .B(_02362_),
    .C(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__a21o_1 _08153_ (.A1(_02361_),
    .A2(_02362_),
    .B1(_02363_),
    .X(_02365_));
 sky130_fd_sc_hd__a22o_1 _08154_ (.A1(net786),
    .A2(net624),
    .B1(_02364_),
    .B2(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__nand4_2 _08155_ (.A(net786),
    .B(net624),
    .C(_02364_),
    .D(_02365_),
    .Y(_02367_));
 sky130_fd_sc_hd__and3_1 _08156_ (.A(_02351_),
    .B(_02366_),
    .C(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__a21oi_1 _08157_ (.A1(_02366_),
    .A2(_02367_),
    .B1(_02351_),
    .Y(_02369_));
 sky130_fd_sc_hd__a21o_1 _08158_ (.A1(_02366_),
    .A2(_02367_),
    .B1(_02351_),
    .X(_02370_));
 sky130_fd_sc_hd__or3b_1 _08159_ (.A(_02368_),
    .B(_02369_),
    .C_N(_02302_),
    .X(_02371_));
 sky130_fd_sc_hd__o21bai_1 _08160_ (.A1(_02368_),
    .A2(_02369_),
    .B1_N(_02302_),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(_02298_),
    .B(_02301_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand3_2 _08162_ (.A(_02371_),
    .B(_02372_),
    .C(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__a21o_1 _08163_ (.A1(_02371_),
    .A2(_02372_),
    .B1(_02373_),
    .X(_02375_));
 sky130_fd_sc_hd__nand3_1 _08164_ (.A(_02305_),
    .B(_02374_),
    .C(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _08165_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02305_),
    .X(_02377_));
 sky130_fd_sc_hd__o21bai_2 _08166_ (.A1(_02309_),
    .A2(_02311_),
    .B1_N(_02308_),
    .Y(_02378_));
 sky130_fd_sc_hd__a21oi_1 _08167_ (.A1(_02376_),
    .A2(_02377_),
    .B1(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__a311o_1 _08168_ (.A1(_02376_),
    .A2(_02377_),
    .A3(_02378_),
    .B1(_02379_),
    .C1(_02240_),
    .X(_02380_));
 sky130_fd_sc_hd__and2b_1 _08169_ (.A_N(_01846_),
    .B(_01851_),
    .X(_02381_));
 sky130_fd_sc_hd__a311o_1 _08170_ (.A1(_01847_),
    .A2(_01853_),
    .A3(_02243_),
    .B1(_02381_),
    .C1(_01845_),
    .X(_02382_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(_01929_),
    .B(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__or2_1 _08172_ (.A(_01929_),
    .B(_02382_),
    .X(_02384_));
 sky130_fd_sc_hd__a32o_1 _08173_ (.A1(net467),
    .A2(_02383_),
    .A3(_02384_),
    .B1(net485),
    .B2(net3656),
    .X(_02385_));
 sky130_fd_sc_hd__and2b_4 _08174_ (.A_N(_02385_),
    .B(_02380_),
    .X(_02386_));
 sky130_fd_sc_hd__inv_2 _08175_ (.A(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__a21oi_2 _08176_ (.A1(net392),
    .A2(_02387_),
    .B1(_02348_),
    .Y(_02388_));
 sky130_fd_sc_hd__o21a_1 _08177_ (.A1(_02318_),
    .A2(_02319_),
    .B1(_02320_),
    .X(_02389_));
 sky130_fd_sc_hd__nor2_1 _08178_ (.A(net3452),
    .B(net3297),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_1 _08179_ (.A(net3452),
    .B(net3297),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2b_1 _08180_ (.A_N(_02390_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__xnor2_1 _08181_ (.A(_02389_),
    .B(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__a21oi_1 _08182_ (.A1(net3582),
    .A2(net403),
    .B1(net362),
    .Y(_02394_));
 sky130_fd_sc_hd__o221a_1 _08183_ (.A1(net373),
    .A2(_02388_),
    .B1(_02393_),
    .B2(net365),
    .C1(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__a21oi_1 _08184_ (.A1(net361),
    .A2(_02326_),
    .B1(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__or2_1 _08185_ (.A(net256),
    .B(net442),
    .X(_02397_));
 sky130_fd_sc_hd__o211a_1 _08186_ (.A1(net449),
    .A2(net3583),
    .B1(_02397_),
    .C1(net845),
    .X(_00642_));
 sky130_fd_sc_hd__mux4_1 _08187_ (.A0(\dpath.RF.R[0][7] ),
    .A1(\dpath.RF.R[1][7] ),
    .A2(\dpath.RF.R[2][7] ),
    .A3(\dpath.RF.R[3][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02398_));
 sky130_fd_sc_hd__mux4_1 _08188_ (.A0(\dpath.RF.R[4][7] ),
    .A1(\dpath.RF.R[5][7] ),
    .A2(\dpath.RF.R[6][7] ),
    .A3(\dpath.RF.R[7][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02399_));
 sky130_fd_sc_hd__o21a_1 _08189_ (.A1(net508),
    .A2(_02399_),
    .B1(net506),
    .X(_02400_));
 sky130_fd_sc_hd__o21ai_1 _08190_ (.A1(net529),
    .A2(_02398_),
    .B1(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__mux4_1 _08191_ (.A0(\dpath.RF.R[12][7] ),
    .A1(\dpath.RF.R[13][7] ),
    .A2(\dpath.RF.R[14][7] ),
    .A3(\dpath.RF.R[15][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02402_));
 sky130_fd_sc_hd__mux4_1 _08192_ (.A0(\dpath.RF.R[8][7] ),
    .A1(\dpath.RF.R[9][7] ),
    .A2(\dpath.RF.R[10][7] ),
    .A3(\dpath.RF.R[11][7] ),
    .S0(net561),
    .S1(net542),
    .X(_02403_));
 sky130_fd_sc_hd__or2_1 _08193_ (.A(net529),
    .B(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__o211a_1 _08194_ (.A1(net508),
    .A2(_02402_),
    .B1(_02404_),
    .C1(net521),
    .X(_02405_));
 sky130_fd_sc_hd__nor2_1 _08195_ (.A(net517),
    .B(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__mux4_1 _08196_ (.A0(\dpath.RF.R[16][7] ),
    .A1(\dpath.RF.R[17][7] ),
    .A2(\dpath.RF.R[18][7] ),
    .A3(\dpath.RF.R[19][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02407_));
 sky130_fd_sc_hd__nor2_1 _08197_ (.A(net529),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__mux4_1 _08198_ (.A0(\dpath.RF.R[20][7] ),
    .A1(\dpath.RF.R[21][7] ),
    .A2(\dpath.RF.R[22][7] ),
    .A3(\dpath.RF.R[23][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02409_));
 sky130_fd_sc_hd__nor2_1 _08199_ (.A(net508),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__mux4_1 _08200_ (.A0(\dpath.RF.R[28][7] ),
    .A1(\dpath.RF.R[29][7] ),
    .A2(\dpath.RF.R[30][7] ),
    .A3(\dpath.RF.R[31][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02411_));
 sky130_fd_sc_hd__nor2_1 _08201_ (.A(net508),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__mux4_1 _08202_ (.A0(\dpath.RF.R[24][7] ),
    .A1(\dpath.RF.R[25][7] ),
    .A2(\dpath.RF.R[26][7] ),
    .A3(\dpath.RF.R[27][7] ),
    .S0(net557),
    .S1(net538),
    .X(_02413_));
 sky130_fd_sc_hd__o21ai_1 _08203_ (.A1(net529),
    .A2(_02413_),
    .B1(net521),
    .Y(_02414_));
 sky130_fd_sc_hd__o32a_1 _08204_ (.A1(net521),
    .A2(_02408_),
    .A3(_02410_),
    .B1(_02412_),
    .B2(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__a221o_1 _08205_ (.A1(_02401_),
    .A2(_02406_),
    .B1(_02415_),
    .B2(net517),
    .C1(net482),
    .X(_02416_));
 sky130_fd_sc_hd__nor2_1 _08206_ (.A(net372),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__mux2_1 _08207_ (.A0(net3654),
    .A1(net30),
    .S(net480),
    .X(_02418_));
 sky130_fd_sc_hd__a221o_1 _08208_ (.A1(net704),
    .A2(net370),
    .B1(net368),
    .B2(_02418_),
    .C1(_02417_),
    .X(_02419_));
 sky130_fd_sc_hd__nand2_1 _08209_ (.A(_02364_),
    .B(_02367_),
    .Y(_02420_));
 sky130_fd_sc_hd__nand4_2 _08210_ (.A(net650),
    .B(net646),
    .C(net765),
    .D(net762),
    .Y(_02421_));
 sky130_fd_sc_hd__a22o_1 _08211_ (.A1(net646),
    .A2(net765),
    .B1(net762),
    .B2(net650),
    .X(_02422_));
 sky130_fd_sc_hd__nand4_2 _08212_ (.A(net641),
    .B(net770),
    .C(_02421_),
    .D(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__a22o_1 _08213_ (.A1(net641),
    .A2(net770),
    .B1(_02421_),
    .B2(_02422_),
    .X(_02424_));
 sky130_fd_sc_hd__and3_1 _08214_ (.A(_02350_),
    .B(_02423_),
    .C(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__inv_2 _08215_ (.A(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__a21oi_1 _08216_ (.A1(_02423_),
    .A2(_02424_),
    .B1(_02350_),
    .Y(_02427_));
 sky130_fd_sc_hd__or2_1 _08217_ (.A(_02425_),
    .B(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__o21bai_1 _08218_ (.A1(_02352_),
    .A2(_02360_),
    .B1_N(_02359_),
    .Y(_02429_));
 sky130_fd_sc_hd__and2_1 _08219_ (.A(net781),
    .B(net628),
    .X(_02430_));
 sky130_fd_sc_hd__nand4_2 _08220_ (.A(net636),
    .B(net776),
    .C(net632),
    .D(net772),
    .Y(_02431_));
 sky130_fd_sc_hd__a22o_1 _08221_ (.A1(net776),
    .A2(net632),
    .B1(net772),
    .B2(net636),
    .X(_02432_));
 sky130_fd_sc_hd__nand3_1 _08222_ (.A(_02430_),
    .B(_02431_),
    .C(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__a21o_1 _08223_ (.A1(_02431_),
    .A2(_02432_),
    .B1(_02430_),
    .X(_02434_));
 sky130_fd_sc_hd__a21bo_1 _08224_ (.A1(_02353_),
    .A2(_02355_),
    .B1_N(_02354_),
    .X(_02435_));
 sky130_fd_sc_hd__and3_1 _08225_ (.A(_02433_),
    .B(_02434_),
    .C(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__nand3_1 _08226_ (.A(_02433_),
    .B(_02434_),
    .C(_02435_),
    .Y(_02437_));
 sky130_fd_sc_hd__a21o_1 _08227_ (.A1(_02433_),
    .A2(_02434_),
    .B1(_02435_),
    .X(_02438_));
 sky130_fd_sc_hd__nand4_1 _08228_ (.A(net783),
    .B(net624),
    .C(_02437_),
    .D(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__a22o_1 _08229_ (.A1(net783),
    .A2(net624),
    .B1(_02437_),
    .B2(_02438_),
    .X(_02440_));
 sky130_fd_sc_hd__and3_1 _08230_ (.A(_02429_),
    .B(_02439_),
    .C(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__a21oi_1 _08231_ (.A1(_02439_),
    .A2(_02440_),
    .B1(_02429_),
    .Y(_02442_));
 sky130_fd_sc_hd__nor2_1 _08232_ (.A(_02441_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(net786),
    .B(net620),
    .Y(_02444_));
 sky130_fd_sc_hd__xor2_2 _08234_ (.A(_02443_),
    .B(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__xor2_1 _08235_ (.A(_02428_),
    .B(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__a21oi_1 _08236_ (.A1(_02302_),
    .A2(_02370_),
    .B1(_02368_),
    .Y(_02447_));
 sky130_fd_sc_hd__xnor2_1 _08237_ (.A(_02446_),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand2_1 _08238_ (.A(_02420_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__xnor2_1 _08239_ (.A(_02420_),
    .B(_02448_),
    .Y(_02450_));
 sky130_fd_sc_hd__xnor2_1 _08240_ (.A(_02374_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__a21bo_1 _08241_ (.A1(_02377_),
    .A2(_02378_),
    .B1_N(_02376_),
    .X(_02452_));
 sky130_fd_sc_hd__and2b_1 _08242_ (.A_N(_02451_),
    .B(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__and2b_1 _08243_ (.A_N(_02452_),
    .B(_02451_),
    .X(_02454_));
 sky130_fd_sc_hd__and3_1 _08244_ (.A(_01926_),
    .B(_01935_),
    .C(_02383_),
    .X(_02455_));
 sky130_fd_sc_hd__a21oi_1 _08245_ (.A1(_01926_),
    .A2(_02383_),
    .B1(_01935_),
    .Y(_02456_));
 sky130_fd_sc_hd__o32a_1 _08246_ (.A1(_02240_),
    .A2(_02453_),
    .A3(_02454_),
    .B1(net484),
    .B2(_01785_),
    .X(_02457_));
 sky130_fd_sc_hd__o31a_4 _08247_ (.A1(net468),
    .A2(_02455_),
    .A3(_02456_),
    .B1(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__inv_2 _08248_ (.A(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__a21oi_4 _08249_ (.A1(net392),
    .A2(_02459_),
    .B1(_02419_),
    .Y(_02460_));
 sky130_fd_sc_hd__nor2_1 _08250_ (.A(net373),
    .B(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__o21a_1 _08251_ (.A1(_02389_),
    .A2(_02390_),
    .B1(_02391_),
    .X(_02462_));
 sky130_fd_sc_hd__nor2_1 _08252_ (.A(net3420),
    .B(net3277),
    .Y(_02463_));
 sky130_fd_sc_hd__nand2_1 _08253_ (.A(net3420),
    .B(net3277),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2b_1 _08254_ (.A_N(_02463_),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__xnor2_1 _08255_ (.A(_02462_),
    .B(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__nor2_1 _08256_ (.A(net365),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__and3_1 _08257_ (.A(net3514),
    .B(net256),
    .C(_02261_),
    .X(_02468_));
 sky130_fd_sc_hd__inv_2 _08258_ (.A(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__a31o_1 _08259_ (.A1(net256),
    .A2(net3280),
    .A3(_02256_),
    .B1(net3514),
    .X(_02470_));
 sky130_fd_sc_hd__a32o_1 _08260_ (.A1(net361),
    .A2(_02469_),
    .A3(_02470_),
    .B1(net403),
    .B2(\dpath.btarg_DX.q[7] ),
    .X(_02471_));
 sky130_fd_sc_hd__or3_1 _08261_ (.A(net450),
    .B(_02467_),
    .C(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__o221a_1 _08262_ (.A1(net3514),
    .A2(net442),
    .B1(_02461_),
    .B2(_02472_),
    .C1(net845),
    .X(_00643_));
 sky130_fd_sc_hd__and2_1 _08263_ (.A(net3473),
    .B(_02468_),
    .X(_02473_));
 sky130_fd_sc_hd__nor2_1 _08264_ (.A(net3473),
    .B(_02468_),
    .Y(_02474_));
 sky130_fd_sc_hd__o21a_1 _08265_ (.A1(_02473_),
    .A2(_02474_),
    .B1(net361),
    .X(_02475_));
 sky130_fd_sc_hd__mux4_1 _08266_ (.A0(\dpath.RF.R[0][8] ),
    .A1(\dpath.RF.R[1][8] ),
    .A2(\dpath.RF.R[2][8] ),
    .A3(\dpath.RF.R[3][8] ),
    .S0(net564),
    .S1(net545),
    .X(_02476_));
 sky130_fd_sc_hd__mux4_1 _08267_ (.A0(\dpath.RF.R[4][8] ),
    .A1(\dpath.RF.R[5][8] ),
    .A2(\dpath.RF.R[6][8] ),
    .A3(\dpath.RF.R[7][8] ),
    .S0(net564),
    .S1(net545),
    .X(_02477_));
 sky130_fd_sc_hd__o21a_1 _08268_ (.A1(net512),
    .A2(_02477_),
    .B1(net506),
    .X(_02478_));
 sky130_fd_sc_hd__o21ai_1 _08269_ (.A1(net532),
    .A2(_02476_),
    .B1(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__mux4_1 _08270_ (.A0(\dpath.RF.R[12][8] ),
    .A1(\dpath.RF.R[13][8] ),
    .A2(\dpath.RF.R[14][8] ),
    .A3(\dpath.RF.R[15][8] ),
    .S0(net564),
    .S1(net545),
    .X(_02480_));
 sky130_fd_sc_hd__mux4_1 _08271_ (.A0(\dpath.RF.R[8][8] ),
    .A1(\dpath.RF.R[9][8] ),
    .A2(\dpath.RF.R[10][8] ),
    .A3(\dpath.RF.R[11][8] ),
    .S0(net565),
    .S1(net544),
    .X(_02481_));
 sky130_fd_sc_hd__or2_1 _08272_ (.A(net532),
    .B(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__o211a_1 _08273_ (.A1(net511),
    .A2(_02480_),
    .B1(_02482_),
    .C1(net523),
    .X(_02483_));
 sky130_fd_sc_hd__nor2_1 _08274_ (.A(net518),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__mux4_1 _08275_ (.A0(\dpath.RF.R[16][8] ),
    .A1(\dpath.RF.R[17][8] ),
    .A2(\dpath.RF.R[18][8] ),
    .A3(\dpath.RF.R[19][8] ),
    .S0(net576),
    .S1(net545),
    .X(_02485_));
 sky130_fd_sc_hd__nor2_1 _08276_ (.A(net532),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__mux4_1 _08277_ (.A0(\dpath.RF.R[20][8] ),
    .A1(\dpath.RF.R[21][8] ),
    .A2(\dpath.RF.R[22][8] ),
    .A3(\dpath.RF.R[23][8] ),
    .S0(net564),
    .S1(net545),
    .X(_02487_));
 sky130_fd_sc_hd__nor2_1 _08278_ (.A(net512),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__mux4_1 _08279_ (.A0(\dpath.RF.R[28][8] ),
    .A1(\dpath.RF.R[29][8] ),
    .A2(\dpath.RF.R[30][8] ),
    .A3(\dpath.RF.R[31][8] ),
    .S0(net564),
    .S1(net545),
    .X(_02489_));
 sky130_fd_sc_hd__nor2_1 _08280_ (.A(net512),
    .B(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__mux4_1 _08281_ (.A0(\dpath.RF.R[24][8] ),
    .A1(\dpath.RF.R[25][8] ),
    .A2(\dpath.RF.R[26][8] ),
    .A3(\dpath.RF.R[27][8] ),
    .S0(net564),
    .S1(net545),
    .X(_02491_));
 sky130_fd_sc_hd__o21ai_1 _08282_ (.A1(net532),
    .A2(_02491_),
    .B1(net524),
    .Y(_02492_));
 sky130_fd_sc_hd__o32a_1 _08283_ (.A1(net524),
    .A2(_02486_),
    .A3(_02488_),
    .B1(_02490_),
    .B2(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__a221o_1 _08284_ (.A1(_02479_),
    .A2(_02484_),
    .B1(_02493_),
    .B2(net518),
    .C1(net482),
    .X(_02494_));
 sky130_fd_sc_hd__nor2_1 _08285_ (.A(net372),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__mux2_2 _08286_ (.A0(net3645),
    .A1(net31),
    .S(net480),
    .X(_02496_));
 sky130_fd_sc_hd__a221o_1 _08287_ (.A1(net703),
    .A2(net370),
    .B1(net368),
    .B2(_02496_),
    .C1(_02495_),
    .X(_02497_));
 sky130_fd_sc_hd__a31o_1 _08288_ (.A1(net786),
    .A2(net620),
    .A3(_02443_),
    .B1(_02441_),
    .X(_02498_));
 sky130_fd_sc_hd__and2_1 _08289_ (.A(_02368_),
    .B(_02446_),
    .X(_02499_));
 sky130_fd_sc_hd__and2_1 _08290_ (.A(net650),
    .B(net757),
    .X(_02500_));
 sky130_fd_sc_hd__and4_1 _08291_ (.A(net646),
    .B(net641),
    .C(net767),
    .D(net762),
    .X(_02501_));
 sky130_fd_sc_hd__nand4_1 _08292_ (.A(net646),
    .B(net641),
    .C(net765),
    .D(net762),
    .Y(_02502_));
 sky130_fd_sc_hd__a22o_1 _08293_ (.A1(net641),
    .A2(net765),
    .B1(net762),
    .B2(net646),
    .X(_02503_));
 sky130_fd_sc_hd__and4_1 _08294_ (.A(net636),
    .B(net770),
    .C(_02502_),
    .D(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__a22o_1 _08295_ (.A1(net636),
    .A2(net770),
    .B1(_02502_),
    .B2(_02503_),
    .X(_02505_));
 sky130_fd_sc_hd__and2b_1 _08296_ (.A_N(_02504_),
    .B(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__nand2_1 _08297_ (.A(_02421_),
    .B(_02423_),
    .Y(_02507_));
 sky130_fd_sc_hd__and2_1 _08298_ (.A(_02506_),
    .B(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__nor2_1 _08299_ (.A(_02506_),
    .B(_02507_),
    .Y(_02509_));
 sky130_fd_sc_hd__or2_1 _08300_ (.A(_02508_),
    .B(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__xnor2_1 _08301_ (.A(_02425_),
    .B(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__a31o_1 _08302_ (.A1(net783),
    .A2(net624),
    .A3(_02438_),
    .B1(_02436_),
    .X(_02512_));
 sky130_fd_sc_hd__and2_1 _08303_ (.A(net781),
    .B(net624),
    .X(_02513_));
 sky130_fd_sc_hd__a22o_1 _08304_ (.A1(net632),
    .A2(net774),
    .B1(net628),
    .B2(net776),
    .X(_02514_));
 sky130_fd_sc_hd__nand4_2 _08305_ (.A(net776),
    .B(net632),
    .C(net774),
    .D(net628),
    .Y(_02515_));
 sky130_fd_sc_hd__nand3_1 _08306_ (.A(_02513_),
    .B(_02514_),
    .C(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__a21o_1 _08307_ (.A1(_02514_),
    .A2(_02515_),
    .B1(_02513_),
    .X(_02517_));
 sky130_fd_sc_hd__a21bo_1 _08308_ (.A1(_02430_),
    .A2(_02432_),
    .B1_N(_02431_),
    .X(_02518_));
 sky130_fd_sc_hd__and3_1 _08309_ (.A(_02516_),
    .B(_02517_),
    .C(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__nand3_1 _08310_ (.A(_02516_),
    .B(_02517_),
    .C(_02518_),
    .Y(_02520_));
 sky130_fd_sc_hd__a21o_1 _08311_ (.A1(_02516_),
    .A2(_02517_),
    .B1(_02518_),
    .X(_02521_));
 sky130_fd_sc_hd__nand4_1 _08312_ (.A(net783),
    .B(net620),
    .C(_02520_),
    .D(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__a22o_1 _08313_ (.A1(net784),
    .A2(net620),
    .B1(_02520_),
    .B2(_02521_),
    .X(_02523_));
 sky130_fd_sc_hd__nand3_2 _08314_ (.A(_02512_),
    .B(_02522_),
    .C(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__a21o_1 _08315_ (.A1(_02522_),
    .A2(_02523_),
    .B1(_02512_),
    .X(_02525_));
 sky130_fd_sc_hd__a22o_1 _08316_ (.A1(net788),
    .A2(net617),
    .B1(_02524_),
    .B2(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__nand4_2 _08317_ (.A(net788),
    .B(net617),
    .C(_02524_),
    .D(_02525_),
    .Y(_02527_));
 sky130_fd_sc_hd__and3_1 _08318_ (.A(_02511_),
    .B(_02526_),
    .C(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__a21oi_1 _08319_ (.A1(_02526_),
    .A2(_02527_),
    .B1(_02511_),
    .Y(_02529_));
 sky130_fd_sc_hd__or4_1 _08320_ (.A(_02428_),
    .B(_02445_),
    .C(_02528_),
    .D(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__o22ai_2 _08321_ (.A1(_02428_),
    .A2(_02445_),
    .B1(_02528_),
    .B2(_02529_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand3_1 _08322_ (.A(_02500_),
    .B(_02530_),
    .C(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__a21o_1 _08323_ (.A1(_02530_),
    .A2(_02531_),
    .B1(_02500_),
    .X(_02533_));
 sky130_fd_sc_hd__and3_1 _08324_ (.A(_02499_),
    .B(_02532_),
    .C(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__a21oi_1 _08325_ (.A1(_02532_),
    .A2(_02533_),
    .B1(_02499_),
    .Y(_02535_));
 sky130_fd_sc_hd__nand2b_1 _08326_ (.A_N(_02371_),
    .B(_02446_),
    .Y(_02536_));
 sky130_fd_sc_hd__or3_1 _08327_ (.A(_02534_),
    .B(_02535_),
    .C(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__o21ai_1 _08328_ (.A1(_02534_),
    .A2(_02535_),
    .B1(_02536_),
    .Y(_02538_));
 sky130_fd_sc_hd__and3_1 _08329_ (.A(_02498_),
    .B(_02537_),
    .C(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__a21oi_1 _08330_ (.A1(_02537_),
    .A2(_02538_),
    .B1(_02498_),
    .Y(_02540_));
 sky130_fd_sc_hd__nor3_1 _08331_ (.A(_02449_),
    .B(_02539_),
    .C(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__o21ai_2 _08332_ (.A1(_02539_),
    .A2(_02540_),
    .B1(_02449_),
    .Y(_02542_));
 sky130_fd_sc_hd__inv_2 _08333_ (.A(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__o21bai_1 _08334_ (.A1(_02374_),
    .A2(_02450_),
    .B1_N(_02453_),
    .Y(_02544_));
 sky130_fd_sc_hd__and3b_1 _08335_ (.A_N(_02541_),
    .B(_02542_),
    .C(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__o21ba_1 _08336_ (.A1(_02541_),
    .A2(_02543_),
    .B1_N(_02544_),
    .X(_02546_));
 sky130_fd_sc_hd__nor3_1 _08337_ (.A(_02240_),
    .B(_02545_),
    .C(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__and3_1 _08338_ (.A(net624),
    .B(net764),
    .C(_01934_),
    .X(_02548_));
 sky130_fd_sc_hd__a311o_1 _08339_ (.A1(_01929_),
    .A2(_01934_),
    .A3(_02382_),
    .B1(_02548_),
    .C1(_01933_),
    .X(_02549_));
 sky130_fd_sc_hd__xnor2_1 _08340_ (.A(_01866_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__a221o_4 _08341_ (.A1(net3416),
    .A2(net485),
    .B1(net467),
    .B2(_02550_),
    .C1(_02547_),
    .X(_02551_));
 sky130_fd_sc_hd__a21oi_4 _08342_ (.A1(net392),
    .A2(_02551_),
    .B1(_02497_),
    .Y(_02552_));
 sky130_fd_sc_hd__o21a_1 _08343_ (.A1(_02462_),
    .A2(_02463_),
    .B1(_02464_),
    .X(_02553_));
 sky130_fd_sc_hd__nor2_1 _08344_ (.A(net3421),
    .B(net3286),
    .Y(_02554_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(net3421),
    .B(net3286),
    .Y(_02555_));
 sky130_fd_sc_hd__nand2b_1 _08346_ (.A_N(_02554_),
    .B(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__xnor2_1 _08347_ (.A(_02553_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__a21oi_1 _08348_ (.A1(\dpath.btarg_DX.q[8] ),
    .A2(_01952_),
    .B1(net362),
    .Y(_02558_));
 sky130_fd_sc_hd__o221a_1 _08349_ (.A1(net373),
    .A2(_02552_),
    .B1(_02557_),
    .B2(net365),
    .C1(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__o21ai_1 _08350_ (.A1(_02475_),
    .A2(_02559_),
    .B1(net442),
    .Y(_02560_));
 sky130_fd_sc_hd__o211a_1 _08351_ (.A1(net3473),
    .A2(net442),
    .B1(_02560_),
    .C1(net845),
    .X(_00644_));
 sky130_fd_sc_hd__and3_1 _08352_ (.A(net3375),
    .B(net3473),
    .C(_02468_),
    .X(_02561_));
 sky130_fd_sc_hd__nor2_1 _08353_ (.A(net3375),
    .B(_02473_),
    .Y(_02562_));
 sky130_fd_sc_hd__o21a_1 _08354_ (.A1(_02561_),
    .A2(_02562_),
    .B1(net361),
    .X(_02563_));
 sky130_fd_sc_hd__mux4_1 _08355_ (.A0(\dpath.RF.R[0][9] ),
    .A1(\dpath.RF.R[1][9] ),
    .A2(\dpath.RF.R[2][9] ),
    .A3(\dpath.RF.R[3][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02564_));
 sky130_fd_sc_hd__mux4_1 _08356_ (.A0(\dpath.RF.R[4][9] ),
    .A1(\dpath.RF.R[5][9] ),
    .A2(\dpath.RF.R[6][9] ),
    .A3(\dpath.RF.R[7][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02565_));
 sky130_fd_sc_hd__o21a_1 _08357_ (.A1(net512),
    .A2(_02565_),
    .B1(net506),
    .X(_02566_));
 sky130_fd_sc_hd__o21ai_1 _08358_ (.A1(net532),
    .A2(_02564_),
    .B1(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__mux4_1 _08359_ (.A0(\dpath.RF.R[12][9] ),
    .A1(\dpath.RF.R[13][9] ),
    .A2(\dpath.RF.R[14][9] ),
    .A3(\dpath.RF.R[15][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02568_));
 sky130_fd_sc_hd__mux4_1 _08360_ (.A0(\dpath.RF.R[8][9] ),
    .A1(\dpath.RF.R[9][9] ),
    .A2(\dpath.RF.R[10][9] ),
    .A3(\dpath.RF.R[11][9] ),
    .S0(net560),
    .S1(net541),
    .X(_02569_));
 sky130_fd_sc_hd__or2_1 _08361_ (.A(net532),
    .B(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__o211a_1 _08362_ (.A1(net511),
    .A2(_02568_),
    .B1(_02570_),
    .C1(net523),
    .X(_02571_));
 sky130_fd_sc_hd__nor2_1 _08363_ (.A(net518),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__mux4_1 _08364_ (.A0(\dpath.RF.R[16][9] ),
    .A1(\dpath.RF.R[17][9] ),
    .A2(\dpath.RF.R[18][9] ),
    .A3(\dpath.RF.R[19][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02573_));
 sky130_fd_sc_hd__nor2_1 _08365_ (.A(net532),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__mux4_1 _08366_ (.A0(\dpath.RF.R[20][9] ),
    .A1(\dpath.RF.R[21][9] ),
    .A2(\dpath.RF.R[22][9] ),
    .A3(\dpath.RF.R[23][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02575_));
 sky130_fd_sc_hd__nor2_1 _08367_ (.A(net512),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__mux4_1 _08368_ (.A0(\dpath.RF.R[28][9] ),
    .A1(\dpath.RF.R[29][9] ),
    .A2(\dpath.RF.R[30][9] ),
    .A3(\dpath.RF.R[31][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02577_));
 sky130_fd_sc_hd__nor2_1 _08369_ (.A(net512),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__mux4_1 _08370_ (.A0(\dpath.RF.R[24][9] ),
    .A1(\dpath.RF.R[25][9] ),
    .A2(\dpath.RF.R[26][9] ),
    .A3(\dpath.RF.R[27][9] ),
    .S0(net565),
    .S1(net544),
    .X(_02579_));
 sky130_fd_sc_hd__o21ai_1 _08371_ (.A1(net532),
    .A2(_02579_),
    .B1(net523),
    .Y(_02580_));
 sky130_fd_sc_hd__o32a_1 _08372_ (.A1(net523),
    .A2(_02574_),
    .A3(_02576_),
    .B1(_02578_),
    .B2(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__a221o_1 _08373_ (.A1(_02567_),
    .A2(_02572_),
    .B1(_02581_),
    .B2(net518),
    .C1(net482),
    .X(_02582_));
 sky130_fd_sc_hd__nor2_1 _08374_ (.A(net372),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__mux2_2 _08375_ (.A0(net3640),
    .A1(net32),
    .S(net480),
    .X(_02584_));
 sky130_fd_sc_hd__a221o_1 _08376_ (.A1(net700),
    .A2(net370),
    .B1(net368),
    .B2(_02584_),
    .C1(_02583_),
    .X(_02585_));
 sky130_fd_sc_hd__a21boi_1 _08377_ (.A1(_01865_),
    .A2(_02549_),
    .B1_N(_01864_),
    .Y(_02586_));
 sky130_fd_sc_hd__or2_1 _08378_ (.A(_01872_),
    .B(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__a21oi_1 _08379_ (.A1(_01872_),
    .A2(_02586_),
    .B1(net468),
    .Y(_02588_));
 sky130_fd_sc_hd__nor2_1 _08380_ (.A(_02541_),
    .B(_02545_),
    .Y(_02589_));
 sky130_fd_sc_hd__a22oi_1 _08381_ (.A1(net646),
    .A2(net757),
    .B1(net754),
    .B2(net650),
    .Y(_02590_));
 sky130_fd_sc_hd__and3_1 _08382_ (.A(net650),
    .B(net646),
    .C(net754),
    .X(_02591_));
 sky130_fd_sc_hd__and2_1 _08383_ (.A(net757),
    .B(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__nor2_1 _08384_ (.A(_02590_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__a31o_1 _08385_ (.A1(net783),
    .A2(net620),
    .A3(_02521_),
    .B1(_02519_),
    .X(_02594_));
 sky130_fd_sc_hd__and2_1 _08386_ (.A(net781),
    .B(net620),
    .X(_02595_));
 sky130_fd_sc_hd__nand4_1 _08387_ (.A(net779),
    .B(net774),
    .C(net628),
    .D(net624),
    .Y(_02596_));
 sky130_fd_sc_hd__a22o_1 _08388_ (.A1(net774),
    .A2(net628),
    .B1(net624),
    .B2(net779),
    .X(_02597_));
 sky130_fd_sc_hd__nand3_1 _08389_ (.A(_02595_),
    .B(_02596_),
    .C(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__a21o_1 _08390_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02595_),
    .X(_02599_));
 sky130_fd_sc_hd__a21bo_1 _08391_ (.A1(_02513_),
    .A2(_02514_),
    .B1_N(_02515_),
    .X(_02600_));
 sky130_fd_sc_hd__and3_1 _08392_ (.A(_02598_),
    .B(_02599_),
    .C(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__nand3_1 _08393_ (.A(_02598_),
    .B(_02599_),
    .C(_02600_),
    .Y(_02602_));
 sky130_fd_sc_hd__a21o_1 _08394_ (.A1(_02598_),
    .A2(_02599_),
    .B1(_02600_),
    .X(_02603_));
 sky130_fd_sc_hd__nand4_1 _08395_ (.A(net785),
    .B(net617),
    .C(_02602_),
    .D(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__a22o_1 _08396_ (.A1(net785),
    .A2(net617),
    .B1(_02602_),
    .B2(_02603_),
    .X(_02605_));
 sky130_fd_sc_hd__nand3_2 _08397_ (.A(_02594_),
    .B(_02604_),
    .C(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__a21o_1 _08398_ (.A1(_02604_),
    .A2(_02605_),
    .B1(_02594_),
    .X(_02607_));
 sky130_fd_sc_hd__a22o_1 _08399_ (.A1(net788),
    .A2(net613),
    .B1(_02606_),
    .B2(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__nand4_2 _08400_ (.A(net788),
    .B(net613),
    .C(_02606_),
    .D(_02607_),
    .Y(_02609_));
 sky130_fd_sc_hd__nor2_1 _08401_ (.A(_02501_),
    .B(_02504_),
    .Y(_02610_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(net632),
    .B(net770),
    .Y(_02611_));
 sky130_fd_sc_hd__and3_1 _08403_ (.A(net641),
    .B(net636),
    .C(net762),
    .X(_02612_));
 sky130_fd_sc_hd__a22o_1 _08404_ (.A1(net636),
    .A2(net765),
    .B1(net762),
    .B2(net641),
    .X(_02613_));
 sky130_fd_sc_hd__a21bo_1 _08405_ (.A1(net767),
    .A2(_02612_),
    .B1_N(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__xor2_2 _08406_ (.A(_02611_),
    .B(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__nand2b_1 _08407_ (.A_N(_02610_),
    .B(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__xnor2_2 _08408_ (.A(_02610_),
    .B(_02615_),
    .Y(_02617_));
 sky130_fd_sc_hd__o21ba_1 _08409_ (.A1(_02426_),
    .A2(_02509_),
    .B1_N(_02508_),
    .X(_02618_));
 sky130_fd_sc_hd__xnor2_1 _08410_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand3_1 _08411_ (.A(_02608_),
    .B(_02609_),
    .C(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__a21o_1 _08412_ (.A1(_02608_),
    .A2(_02609_),
    .B1(_02619_),
    .X(_02621_));
 sky130_fd_sc_hd__nand3_1 _08413_ (.A(_02528_),
    .B(_02620_),
    .C(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__a21o_1 _08414_ (.A1(_02620_),
    .A2(_02621_),
    .B1(_02528_),
    .X(_02623_));
 sky130_fd_sc_hd__nand3_1 _08415_ (.A(_02593_),
    .B(_02622_),
    .C(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__a21o_1 _08416_ (.A1(_02622_),
    .A2(_02623_),
    .B1(_02593_),
    .X(_02625_));
 sky130_fd_sc_hd__a21bo_1 _08417_ (.A1(_02500_),
    .A2(_02531_),
    .B1_N(_02530_),
    .X(_02626_));
 sky130_fd_sc_hd__nand3_2 _08418_ (.A(_02624_),
    .B(_02625_),
    .C(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__a21o_1 _08419_ (.A1(_02624_),
    .A2(_02625_),
    .B1(_02626_),
    .X(_02628_));
 sky130_fd_sc_hd__and3_1 _08420_ (.A(_02534_),
    .B(_02627_),
    .C(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__a21oi_1 _08421_ (.A1(_02627_),
    .A2(_02628_),
    .B1(_02534_),
    .Y(_02630_));
 sky130_fd_sc_hd__a211oi_2 _08422_ (.A1(_02524_),
    .A2(_02527_),
    .B1(_02629_),
    .C1(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__o211a_1 _08423_ (.A1(_02629_),
    .A2(_02630_),
    .B1(_02524_),
    .C1(_02527_),
    .X(_02632_));
 sky130_fd_sc_hd__a21boi_1 _08424_ (.A1(_02498_),
    .A2(_02538_),
    .B1_N(_02537_),
    .Y(_02633_));
 sky130_fd_sc_hd__o21a_1 _08425_ (.A1(_02631_),
    .A2(_02632_),
    .B1(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__o21ai_1 _08426_ (.A1(_02631_),
    .A2(_02632_),
    .B1(_02633_),
    .Y(_02635_));
 sky130_fd_sc_hd__nor3_1 _08427_ (.A(_02631_),
    .B(_02632_),
    .C(_02633_),
    .Y(_02636_));
 sky130_fd_sc_hd__nor2_1 _08428_ (.A(_02634_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__xnor2_1 _08429_ (.A(_02589_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(net3662),
    .A1(_02638_),
    .S(net484),
    .X(_02639_));
 sky130_fd_sc_hd__a22o_4 _08431_ (.A1(_02587_),
    .A2(_02588_),
    .B1(_02639_),
    .B2(net468),
    .X(_02640_));
 sky130_fd_sc_hd__a21oi_4 _08432_ (.A1(net392),
    .A2(_02640_),
    .B1(_02585_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21a_1 _08433_ (.A1(_02553_),
    .A2(_02554_),
    .B1(_02555_),
    .X(_02642_));
 sky130_fd_sc_hd__nor2_1 _08434_ (.A(net3461),
    .B(net3228),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _08435_ (.A(net3461),
    .B(net3228),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2b_1 _08436_ (.A_N(_02643_),
    .B(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__xnor2_1 _08437_ (.A(_02642_),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__a21oi_1 _08438_ (.A1(net3565),
    .A2(_01952_),
    .B1(net361),
    .Y(_02647_));
 sky130_fd_sc_hd__o221a_1 _08439_ (.A1(net373),
    .A2(_02641_),
    .B1(_02646_),
    .B2(net365),
    .C1(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__nor2_1 _08440_ (.A(_02563_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__or2_1 _08441_ (.A(net3375),
    .B(net442),
    .X(_02650_));
 sky130_fd_sc_hd__o211a_1 _08442_ (.A1(net450),
    .A2(_02649_),
    .B1(_02650_),
    .C1(net845),
    .X(_00645_));
 sky130_fd_sc_hd__and2_1 _08443_ (.A(net3587),
    .B(_02561_),
    .X(_02651_));
 sky130_fd_sc_hd__nor2_1 _08444_ (.A(net3587),
    .B(_02561_),
    .Y(_02652_));
 sky130_fd_sc_hd__o21a_1 _08445_ (.A1(_02651_),
    .A2(_02652_),
    .B1(net361),
    .X(_02653_));
 sky130_fd_sc_hd__mux4_1 _08446_ (.A0(\dpath.RF.R[0][10] ),
    .A1(\dpath.RF.R[1][10] ),
    .A2(\dpath.RF.R[2][10] ),
    .A3(\dpath.RF.R[3][10] ),
    .S0(net564),
    .S1(net544),
    .X(_02654_));
 sky130_fd_sc_hd__mux4_1 _08447_ (.A0(\dpath.RF.R[4][10] ),
    .A1(\dpath.RF.R[5][10] ),
    .A2(\dpath.RF.R[6][10] ),
    .A3(\dpath.RF.R[7][10] ),
    .S0(net565),
    .S1(net544),
    .X(_02655_));
 sky130_fd_sc_hd__o21a_1 _08448_ (.A1(net511),
    .A2(_02655_),
    .B1(net506),
    .X(_02656_));
 sky130_fd_sc_hd__o21ai_1 _08449_ (.A1(net531),
    .A2(_02654_),
    .B1(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__mux4_1 _08450_ (.A0(\dpath.RF.R[12][10] ),
    .A1(\dpath.RF.R[13][10] ),
    .A2(\dpath.RF.R[14][10] ),
    .A3(\dpath.RF.R[15][10] ),
    .S0(net564),
    .S1(net544),
    .X(_02658_));
 sky130_fd_sc_hd__mux4_1 _08451_ (.A0(\dpath.RF.R[8][10] ),
    .A1(\dpath.RF.R[9][10] ),
    .A2(\dpath.RF.R[10][10] ),
    .A3(\dpath.RF.R[11][10] ),
    .S0(net565),
    .S1(net544),
    .X(_02659_));
 sky130_fd_sc_hd__or2_1 _08452_ (.A(net531),
    .B(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__o211a_1 _08453_ (.A1(net511),
    .A2(_02658_),
    .B1(_02660_),
    .C1(net523),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_1 _08454_ (.A(net518),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__mux4_1 _08455_ (.A0(\dpath.RF.R[16][10] ),
    .A1(\dpath.RF.R[17][10] ),
    .A2(\dpath.RF.R[18][10] ),
    .A3(\dpath.RF.R[19][10] ),
    .S0(net564),
    .S1(net545),
    .X(_02663_));
 sky130_fd_sc_hd__nor2_1 _08456_ (.A(net531),
    .B(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__mux4_1 _08457_ (.A0(\dpath.RF.R[20][10] ),
    .A1(\dpath.RF.R[21][10] ),
    .A2(\dpath.RF.R[22][10] ),
    .A3(\dpath.RF.R[23][10] ),
    .S0(net564),
    .S1(net545),
    .X(_02665_));
 sky130_fd_sc_hd__nor2_1 _08458_ (.A(net511),
    .B(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__mux4_1 _08459_ (.A0(\dpath.RF.R[28][10] ),
    .A1(\dpath.RF.R[29][10] ),
    .A2(\dpath.RF.R[30][10] ),
    .A3(\dpath.RF.R[31][10] ),
    .S0(net564),
    .S1(net545),
    .X(_02667_));
 sky130_fd_sc_hd__nor2_1 _08460_ (.A(net511),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__mux4_1 _08461_ (.A0(\dpath.RF.R[24][10] ),
    .A1(\dpath.RF.R[25][10] ),
    .A2(\dpath.RF.R[26][10] ),
    .A3(\dpath.RF.R[27][10] ),
    .S0(net564),
    .S1(net545),
    .X(_02669_));
 sky130_fd_sc_hd__o21ai_1 _08462_ (.A1(net531),
    .A2(_02669_),
    .B1(net524),
    .Y(_02670_));
 sky130_fd_sc_hd__o32a_1 _08463_ (.A1(net524),
    .A2(_02664_),
    .A3(_02666_),
    .B1(_02668_),
    .B2(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__a221o_1 _08464_ (.A1(_02657_),
    .A2(_02662_),
    .B1(_02671_),
    .B2(net518),
    .C1(net482),
    .X(_02672_));
 sky130_fd_sc_hd__nor2_1 _08465_ (.A(net372),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__mux2_2 _08466_ (.A0(net3641),
    .A1(net2),
    .S(net479),
    .X(_02674_));
 sky130_fd_sc_hd__a221o_1 _08467_ (.A1(net698),
    .A2(net370),
    .B1(net368),
    .B2(_02674_),
    .C1(_02673_),
    .X(_02675_));
 sky130_fd_sc_hd__nand2_1 _08468_ (.A(_02606_),
    .B(_02609_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _08469_ (.A(net641),
    .B(net757),
    .Y(_02677_));
 sky130_fd_sc_hd__a22o_1 _08470_ (.A1(net646),
    .A2(net754),
    .B1(net751),
    .B2(net650),
    .X(_02678_));
 sky130_fd_sc_hd__a21bo_1 _08471_ (.A1(net751),
    .A2(_02591_),
    .B1_N(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__xor2_1 _08472_ (.A(_02677_),
    .B(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__or3b_1 _08473_ (.A(_02426_),
    .B(_02510_),
    .C_N(_02617_),
    .X(_02681_));
 sky130_fd_sc_hd__nand2_1 _08474_ (.A(_02620_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__a31o_1 _08475_ (.A1(net785),
    .A2(net617),
    .A3(_02603_),
    .B1(_02601_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _08476_ (.A(net785),
    .B(net613),
    .Y(_02684_));
 sky130_fd_sc_hd__and2_1 _08477_ (.A(net781),
    .B(net617),
    .X(_02685_));
 sky130_fd_sc_hd__a22o_1 _08478_ (.A1(net774),
    .A2(net624),
    .B1(net620),
    .B2(net779),
    .X(_02686_));
 sky130_fd_sc_hd__nand4_1 _08479_ (.A(net779),
    .B(net774),
    .C(net624),
    .D(net620),
    .Y(_02687_));
 sky130_fd_sc_hd__nand3_1 _08480_ (.A(_02685_),
    .B(_02686_),
    .C(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__a21o_1 _08481_ (.A1(_02686_),
    .A2(_02687_),
    .B1(_02685_),
    .X(_02689_));
 sky130_fd_sc_hd__a21bo_1 _08482_ (.A1(_02595_),
    .A2(_02597_),
    .B1_N(_02596_),
    .X(_02690_));
 sky130_fd_sc_hd__nand3_1 _08483_ (.A(_02688_),
    .B(_02689_),
    .C(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21o_1 _08484_ (.A1(_02688_),
    .A2(_02689_),
    .B1(_02690_),
    .X(_02692_));
 sky130_fd_sc_hd__nand3b_2 _08485_ (.A_N(_02684_),
    .B(_02691_),
    .C(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__a21bo_1 _08486_ (.A1(_02691_),
    .A2(_02692_),
    .B1_N(_02684_),
    .X(_02694_));
 sky130_fd_sc_hd__nand3_4 _08487_ (.A(_02683_),
    .B(_02693_),
    .C(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__a21o_1 _08488_ (.A1(_02693_),
    .A2(_02694_),
    .B1(_02683_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_1 _08489_ (.A(net788),
    .B(net611),
    .X(_02697_));
 sky130_fd_sc_hd__a21o_1 _08490_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__nand3_2 _08491_ (.A(_02695_),
    .B(_02696_),
    .C(_02697_),
    .Y(_02699_));
 sky130_fd_sc_hd__and2_1 _08492_ (.A(_02698_),
    .B(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__a32o_1 _08493_ (.A1(net632),
    .A2(net770),
    .A3(_02613_),
    .B1(_02612_),
    .B2(net767),
    .X(_02701_));
 sky130_fd_sc_hd__a22o_1 _08494_ (.A1(net632),
    .A2(net765),
    .B1(net762),
    .B2(net636),
    .X(_02702_));
 sky130_fd_sc_hd__nand4_2 _08495_ (.A(net636),
    .B(net632),
    .C(net765),
    .D(net762),
    .Y(_02703_));
 sky130_fd_sc_hd__nand3_1 _08496_ (.A(_01845_),
    .B(_02702_),
    .C(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__a21o_1 _08497_ (.A1(_02702_),
    .A2(_02703_),
    .B1(_01845_),
    .X(_02705_));
 sky130_fd_sc_hd__nand3_1 _08498_ (.A(_02592_),
    .B(_02704_),
    .C(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__a21o_1 _08499_ (.A1(_02704_),
    .A2(_02705_),
    .B1(_02592_),
    .X(_02707_));
 sky130_fd_sc_hd__and3_1 _08500_ (.A(_02701_),
    .B(_02706_),
    .C(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__a21oi_1 _08501_ (.A1(_02706_),
    .A2(_02707_),
    .B1(_02701_),
    .Y(_02709_));
 sky130_fd_sc_hd__or2_1 _08502_ (.A(_02708_),
    .B(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(_02508_),
    .B(_02617_),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2_1 _08504_ (.A(_02616_),
    .B(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__xnor2_1 _08505_ (.A(_02710_),
    .B(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__nand2_1 _08506_ (.A(_02700_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__xnor2_1 _08507_ (.A(_02700_),
    .B(_02713_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand2b_1 _08508_ (.A_N(_02715_),
    .B(_02682_),
    .Y(_02716_));
 sky130_fd_sc_hd__xnor2_1 _08509_ (.A(_02682_),
    .B(_02715_),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2_1 _08510_ (.A(_02680_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__xor2_1 _08511_ (.A(_02680_),
    .B(_02717_),
    .X(_02719_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(_02622_),
    .B(_02624_),
    .Y(_02720_));
 sky130_fd_sc_hd__nand2_1 _08513_ (.A(_02719_),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__xor2_1 _08514_ (.A(_02719_),
    .B(_02720_),
    .X(_02722_));
 sky130_fd_sc_hd__and2b_1 _08515_ (.A_N(_02627_),
    .B(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__xnor2_1 _08516_ (.A(_02627_),
    .B(_02722_),
    .Y(_02724_));
 sky130_fd_sc_hd__and2_1 _08517_ (.A(_02676_),
    .B(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__xnor2_1 _08518_ (.A(_02676_),
    .B(_02724_),
    .Y(_02726_));
 sky130_fd_sc_hd__or2_1 _08519_ (.A(_02629_),
    .B(_02631_),
    .X(_02727_));
 sky130_fd_sc_hd__and2b_1 _08520_ (.A_N(_02726_),
    .B(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__xor2_1 _08521_ (.A(_02726_),
    .B(_02727_),
    .X(_02729_));
 sky130_fd_sc_hd__a211o_1 _08522_ (.A1(_02542_),
    .A2(_02544_),
    .B1(_02636_),
    .C1(_02541_),
    .X(_02730_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(_02635_),
    .B(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__and3b_1 _08524_ (.A_N(_02729_),
    .B(_02730_),
    .C(_02635_),
    .X(_02732_));
 sky130_fd_sc_hd__a211o_1 _08525_ (.A1(_02729_),
    .A2(_02731_),
    .B1(_02732_),
    .C1(_02240_),
    .X(_02733_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(net3483),
    .B(net485),
    .Y(_02734_));
 sky130_fd_sc_hd__nor2_1 _08527_ (.A(_01864_),
    .B(_01871_),
    .Y(_02735_));
 sky130_fd_sc_hd__and4b_1 _08528_ (.A_N(_01872_),
    .B(_02549_),
    .C(_01864_),
    .D(_01865_),
    .X(_02736_));
 sky130_fd_sc_hd__o31a_1 _08529_ (.A1(_01870_),
    .A2(_02735_),
    .A3(_02736_),
    .B1(_01925_),
    .X(_02737_));
 sky130_fd_sc_hd__nor4_1 _08530_ (.A(_01870_),
    .B(_01925_),
    .C(_02735_),
    .D(_02736_),
    .Y(_02738_));
 sky130_fd_sc_hd__o311a_4 _08531_ (.A1(net468),
    .A2(_02737_),
    .A3(_02738_),
    .B1(_02733_),
    .C1(net3484),
    .X(_02739_));
 sky130_fd_sc_hd__inv_2 _08532_ (.A(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__a21oi_4 _08533_ (.A1(net392),
    .A2(_02740_),
    .B1(_02675_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_1 _08534_ (.A(net3435),
    .B(net3274),
    .Y(_02742_));
 sky130_fd_sc_hd__or2_1 _08535_ (.A(net3435),
    .B(net3274),
    .X(_02743_));
 sky130_fd_sc_hd__nand2_1 _08536_ (.A(_02742_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__o21ai_1 _08537_ (.A1(_02642_),
    .A2(_02643_),
    .B1(_02644_),
    .Y(_02745_));
 sky130_fd_sc_hd__xor2_1 _08538_ (.A(_02744_),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__a21oi_1 _08539_ (.A1(\dpath.btarg_DX.q[10] ),
    .A2(net403),
    .B1(net361),
    .Y(_02747_));
 sky130_fd_sc_hd__o221a_1 _08540_ (.A1(net373),
    .A2(_02741_),
    .B1(_02746_),
    .B2(net365),
    .C1(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__nor2_1 _08541_ (.A(_02653_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__or2_1 _08542_ (.A(net3587),
    .B(net441),
    .X(_02750_));
 sky130_fd_sc_hd__o211a_1 _08543_ (.A1(net449),
    .A2(_02749_),
    .B1(_02750_),
    .C1(net845),
    .X(_00646_));
 sky130_fd_sc_hd__and3_1 _08544_ (.A(net3410),
    .B(net229),
    .C(_02561_),
    .X(_02751_));
 sky130_fd_sc_hd__nor2_1 _08545_ (.A(net3410),
    .B(_02651_),
    .Y(_02752_));
 sky130_fd_sc_hd__o21a_1 _08546_ (.A1(_02751_),
    .A2(_02752_),
    .B1(net361),
    .X(_02753_));
 sky130_fd_sc_hd__mux4_1 _08547_ (.A0(\dpath.RF.R[0][11] ),
    .A1(\dpath.RF.R[1][11] ),
    .A2(\dpath.RF.R[2][11] ),
    .A3(\dpath.RF.R[3][11] ),
    .S0(net561),
    .S1(net542),
    .X(_02754_));
 sky130_fd_sc_hd__mux4_1 _08548_ (.A0(\dpath.RF.R[4][11] ),
    .A1(\dpath.RF.R[5][11] ),
    .A2(\dpath.RF.R[6][11] ),
    .A3(\dpath.RF.R[7][11] ),
    .S0(net557),
    .S1(net538),
    .X(_02755_));
 sky130_fd_sc_hd__o21a_1 _08549_ (.A1(net508),
    .A2(_02755_),
    .B1(net506),
    .X(_02756_));
 sky130_fd_sc_hd__o21ai_1 _08550_ (.A1(net529),
    .A2(_02754_),
    .B1(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__mux4_1 _08551_ (.A0(\dpath.RF.R[12][11] ),
    .A1(\dpath.RF.R[13][11] ),
    .A2(\dpath.RF.R[14][11] ),
    .A3(\dpath.RF.R[15][11] ),
    .S0(net559),
    .S1(net540),
    .X(_02758_));
 sky130_fd_sc_hd__mux4_1 _08552_ (.A0(\dpath.RF.R[8][11] ),
    .A1(\dpath.RF.R[9][11] ),
    .A2(\dpath.RF.R[10][11] ),
    .A3(\dpath.RF.R[11][11] ),
    .S0(net559),
    .S1(net540),
    .X(_02759_));
 sky130_fd_sc_hd__or2_1 _08553_ (.A(net530),
    .B(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__o211a_1 _08554_ (.A1(net509),
    .A2(_02758_),
    .B1(_02760_),
    .C1(net522),
    .X(_02761_));
 sky130_fd_sc_hd__nor2_1 _08555_ (.A(net517),
    .B(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__mux4_1 _08556_ (.A0(\dpath.RF.R[16][11] ),
    .A1(\dpath.RF.R[17][11] ),
    .A2(\dpath.RF.R[18][11] ),
    .A3(\dpath.RF.R[19][11] ),
    .S0(net559),
    .S1(net540),
    .X(_02763_));
 sky130_fd_sc_hd__nor2_1 _08557_ (.A(net530),
    .B(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__mux4_1 _08558_ (.A0(\dpath.RF.R[20][11] ),
    .A1(\dpath.RF.R[21][11] ),
    .A2(\dpath.RF.R[22][11] ),
    .A3(\dpath.RF.R[23][11] ),
    .S0(net559),
    .S1(net540),
    .X(_02765_));
 sky130_fd_sc_hd__nor2_1 _08559_ (.A(net509),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__mux4_1 _08560_ (.A0(\dpath.RF.R[28][11] ),
    .A1(\dpath.RF.R[29][11] ),
    .A2(\dpath.RF.R[30][11] ),
    .A3(\dpath.RF.R[31][11] ),
    .S0(net559),
    .S1(net540),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _08561_ (.A(net509),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__mux4_1 _08562_ (.A0(\dpath.RF.R[24][11] ),
    .A1(\dpath.RF.R[25][11] ),
    .A2(\dpath.RF.R[26][11] ),
    .A3(\dpath.RF.R[27][11] ),
    .S0(net559),
    .S1(net540),
    .X(_02769_));
 sky130_fd_sc_hd__o21ai_1 _08563_ (.A1(net530),
    .A2(_02769_),
    .B1(net521),
    .Y(_02770_));
 sky130_fd_sc_hd__o32a_1 _08564_ (.A1(net521),
    .A2(_02764_),
    .A3(_02766_),
    .B1(_02768_),
    .B2(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__a221o_1 _08565_ (.A1(_02757_),
    .A2(_02762_),
    .B1(_02771_),
    .B2(net517),
    .C1(net482),
    .X(_02772_));
 sky130_fd_sc_hd__nor2_1 _08566_ (.A(net372),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__mux2_1 _08567_ (.A0(net3648),
    .A1(net3),
    .S(net480),
    .X(_02774_));
 sky130_fd_sc_hd__a221o_1 _08568_ (.A1(net3627),
    .A2(net370),
    .B1(net368),
    .B2(_02774_),
    .C1(_02773_),
    .X(_02775_));
 sky130_fd_sc_hd__or3_1 _08569_ (.A(_01887_),
    .B(_01923_),
    .C(_02737_),
    .X(_02776_));
 sky130_fd_sc_hd__o21ai_2 _08570_ (.A1(_01923_),
    .A2(_02737_),
    .B1(_01887_),
    .Y(_02777_));
 sky130_fd_sc_hd__or2_1 _08571_ (.A(_02728_),
    .B(_02732_),
    .X(_02778_));
 sky130_fd_sc_hd__nand2_1 _08572_ (.A(net636),
    .B(net757),
    .Y(_02779_));
 sky130_fd_sc_hd__a22o_1 _08573_ (.A1(net641),
    .A2(net754),
    .B1(net751),
    .B2(net646),
    .X(_02780_));
 sky130_fd_sc_hd__and3_1 _08574_ (.A(net646),
    .B(net641),
    .C(net751),
    .X(_02781_));
 sky130_fd_sc_hd__a21bo_1 _08575_ (.A1(net754),
    .A2(_02781_),
    .B1_N(_02780_),
    .X(_02782_));
 sky130_fd_sc_hd__xor2_1 _08576_ (.A(_02779_),
    .B(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__and3_1 _08577_ (.A(net650),
    .B(net748),
    .C(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__a21oi_1 _08578_ (.A1(net650),
    .A2(net748),
    .B1(_02783_),
    .Y(_02785_));
 sky130_fd_sc_hd__or2_1 _08579_ (.A(_02784_),
    .B(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__or2_1 _08580_ (.A(_02710_),
    .B(_02711_),
    .X(_02787_));
 sky130_fd_sc_hd__nand2_1 _08581_ (.A(_02691_),
    .B(_02693_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _08582_ (.A(net785),
    .B(net611),
    .Y(_02789_));
 sky130_fd_sc_hd__and2_1 _08583_ (.A(net781),
    .B(net613),
    .X(_02790_));
 sky130_fd_sc_hd__a22o_1 _08584_ (.A1(net774),
    .A2(net620),
    .B1(net617),
    .B2(net779),
    .X(_02791_));
 sky130_fd_sc_hd__nand4_2 _08585_ (.A(net779),
    .B(net774),
    .C(net620),
    .D(net617),
    .Y(_02792_));
 sky130_fd_sc_hd__nand3_1 _08586_ (.A(_02790_),
    .B(_02791_),
    .C(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__a21o_1 _08587_ (.A1(_02791_),
    .A2(_02792_),
    .B1(_02790_),
    .X(_02794_));
 sky130_fd_sc_hd__a21bo_1 _08588_ (.A1(_02685_),
    .A2(_02686_),
    .B1_N(_02687_),
    .X(_02795_));
 sky130_fd_sc_hd__and3_1 _08589_ (.A(_02793_),
    .B(_02794_),
    .C(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__a21oi_1 _08590_ (.A1(_02793_),
    .A2(_02794_),
    .B1(_02795_),
    .Y(_02797_));
 sky130_fd_sc_hd__nor2_1 _08591_ (.A(_02796_),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__xnor2_1 _08592_ (.A(_02789_),
    .B(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__and2_1 _08593_ (.A(_02788_),
    .B(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__xor2_1 _08594_ (.A(_02788_),
    .B(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__nand2_1 _08595_ (.A(net788),
    .B(net608),
    .Y(_02802_));
 sky130_fd_sc_hd__and3_1 _08596_ (.A(net789),
    .B(net608),
    .C(_02801_),
    .X(_02803_));
 sky130_fd_sc_hd__xor2_1 _08597_ (.A(_02801_),
    .B(_02802_),
    .X(_02804_));
 sky130_fd_sc_hd__nor2_1 _08598_ (.A(_02616_),
    .B(_02710_),
    .Y(_02805_));
 sky130_fd_sc_hd__a21boi_1 _08599_ (.A1(_02701_),
    .A2(_02707_),
    .B1_N(_02706_),
    .Y(_02806_));
 sky130_fd_sc_hd__nand2_1 _08600_ (.A(_02703_),
    .B(_02704_),
    .Y(_02807_));
 sky130_fd_sc_hd__a32o_1 _08601_ (.A1(net641),
    .A2(net757),
    .A3(_02678_),
    .B1(_02591_),
    .B2(net751),
    .X(_02808_));
 sky130_fd_sc_hd__a22o_1 _08602_ (.A1(net628),
    .A2(net765),
    .B1(net762),
    .B2(net632),
    .X(_02809_));
 sky130_fd_sc_hd__nand4_2 _08603_ (.A(net632),
    .B(net628),
    .C(net765),
    .D(net762),
    .Y(_02810_));
 sky130_fd_sc_hd__nand4_1 _08604_ (.A(net770),
    .B(net624),
    .C(_02809_),
    .D(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__a22o_1 _08605_ (.A1(net770),
    .A2(net624),
    .B1(_02809_),
    .B2(_02810_),
    .X(_02812_));
 sky130_fd_sc_hd__nand2_1 _08606_ (.A(_02811_),
    .B(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__xnor2_1 _08607_ (.A(_02808_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__xor2_1 _08608_ (.A(_02807_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__nand2b_1 _08609_ (.A_N(_02806_),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__xnor2_1 _08610_ (.A(_02806_),
    .B(_02815_),
    .Y(_02817_));
 sky130_fd_sc_hd__nand2_1 _08611_ (.A(_02805_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__xnor2_1 _08612_ (.A(_02805_),
    .B(_02817_),
    .Y(_02819_));
 sky130_fd_sc_hd__or2_1 _08613_ (.A(_02804_),
    .B(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__xnor2_1 _08614_ (.A(_02804_),
    .B(_02819_),
    .Y(_02821_));
 sky130_fd_sc_hd__a21oi_2 _08615_ (.A1(_02714_),
    .A2(_02787_),
    .B1(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__and3_1 _08616_ (.A(_02714_),
    .B(_02787_),
    .C(_02821_),
    .X(_02823_));
 sky130_fd_sc_hd__nor3_2 _08617_ (.A(_02786_),
    .B(_02822_),
    .C(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__o21a_1 _08618_ (.A1(_02822_),
    .A2(_02823_),
    .B1(_02786_),
    .X(_02825_));
 sky130_fd_sc_hd__a211oi_2 _08619_ (.A1(_02716_),
    .A2(_02718_),
    .B1(_02824_),
    .C1(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__o211a_1 _08620_ (.A1(_02824_),
    .A2(_02825_),
    .B1(_02716_),
    .C1(_02718_),
    .X(_02827_));
 sky130_fd_sc_hd__nor3_2 _08621_ (.A(_02721_),
    .B(_02826_),
    .C(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__o21a_1 _08622_ (.A1(_02826_),
    .A2(_02827_),
    .B1(_02721_),
    .X(_02829_));
 sky130_fd_sc_hd__a211oi_2 _08623_ (.A1(_02695_),
    .A2(_02699_),
    .B1(_02828_),
    .C1(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__a211o_1 _08624_ (.A1(_02695_),
    .A2(_02699_),
    .B1(_02828_),
    .C1(_02829_),
    .X(_02831_));
 sky130_fd_sc_hd__o211ai_2 _08625_ (.A1(_02828_),
    .A2(_02829_),
    .B1(_02695_),
    .C1(_02699_),
    .Y(_02832_));
 sky130_fd_sc_hd__a211o_1 _08626_ (.A1(_02831_),
    .A2(_02832_),
    .B1(_02723_),
    .C1(_02725_),
    .X(_02833_));
 sky130_fd_sc_hd__o211a_2 _08627_ (.A1(_02723_),
    .A2(_02725_),
    .B1(_02831_),
    .C1(_02832_),
    .X(_02834_));
 sky130_fd_sc_hd__inv_2 _08628_ (.A(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _08629_ (.A(_02833_),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__xnor2_1 _08630_ (.A(_02778_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__or2_1 _08631_ (.A(net3685),
    .B(net484),
    .X(_02838_));
 sky130_fd_sc_hd__o211a_1 _08632_ (.A1(net485),
    .A2(_02837_),
    .B1(_02838_),
    .C1(net468),
    .X(_02839_));
 sky130_fd_sc_hd__a31o_4 _08633_ (.A1(net467),
    .A2(_02776_),
    .A3(_02777_),
    .B1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__a21oi_4 _08634_ (.A1(net392),
    .A2(_02840_),
    .B1(net3628),
    .Y(_02841_));
 sky130_fd_sc_hd__nor2_4 _08635_ (.A(net481),
    .B(_02126_),
    .Y(_02842_));
 sky130_fd_sc_hd__inv_2 _08636_ (.A(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__nand2_4 _08637_ (.A(net578),
    .B(_02125_),
    .Y(_02844_));
 sky130_fd_sc_hd__a21bo_1 _08638_ (.A1(_02126_),
    .A2(_02128_),
    .B1_N(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__and2_1 _08639_ (.A(net3358),
    .B(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__xor2_1 _08640_ (.A(net3358),
    .B(_02845_),
    .X(_02847_));
 sky130_fd_sc_hd__a21bo_1 _08641_ (.A1(_02743_),
    .A2(_02745_),
    .B1_N(_02742_),
    .X(_02848_));
 sky130_fd_sc_hd__xnor2_1 _08642_ (.A(_02847_),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__o2bb2a_1 _08643_ (.A1_N(net3426),
    .A2_N(_01952_),
    .B1(net365),
    .B2(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__o211a_1 _08644_ (.A1(net373),
    .A2(_02841_),
    .B1(_02850_),
    .C1(_01958_),
    .X(_02851_));
 sky130_fd_sc_hd__o21ai_1 _08645_ (.A1(_02753_),
    .A2(net3427),
    .B1(net441),
    .Y(_02852_));
 sky130_fd_sc_hd__o211a_1 _08646_ (.A1(net3410),
    .A2(net441),
    .B1(net3428),
    .C1(net845),
    .X(_00647_));
 sky130_fd_sc_hd__xnor2_1 _08647_ (.A(net3579),
    .B(_02751_),
    .Y(_02853_));
 sky130_fd_sc_hd__mux4_1 _08648_ (.A0(\dpath.RF.R[0][12] ),
    .A1(\dpath.RF.R[1][12] ),
    .A2(\dpath.RF.R[2][12] ),
    .A3(\dpath.RF.R[3][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02854_));
 sky130_fd_sc_hd__mux4_1 _08649_ (.A0(\dpath.RF.R[4][12] ),
    .A1(\dpath.RF.R[5][12] ),
    .A2(\dpath.RF.R[6][12] ),
    .A3(\dpath.RF.R[7][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02855_));
 sky130_fd_sc_hd__o21a_1 _08650_ (.A1(net509),
    .A2(_02855_),
    .B1(net506),
    .X(_02856_));
 sky130_fd_sc_hd__o21ai_1 _08651_ (.A1(net530),
    .A2(_02854_),
    .B1(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__mux4_1 _08652_ (.A0(\dpath.RF.R[12][12] ),
    .A1(\dpath.RF.R[13][12] ),
    .A2(\dpath.RF.R[14][12] ),
    .A3(\dpath.RF.R[15][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02858_));
 sky130_fd_sc_hd__mux4_1 _08653_ (.A0(\dpath.RF.R[8][12] ),
    .A1(\dpath.RF.R[9][12] ),
    .A2(\dpath.RF.R[10][12] ),
    .A3(\dpath.RF.R[11][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02859_));
 sky130_fd_sc_hd__or2_1 _08654_ (.A(net530),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__o211a_1 _08655_ (.A1(net509),
    .A2(_02858_),
    .B1(_02860_),
    .C1(net522),
    .X(_02861_));
 sky130_fd_sc_hd__nor2_1 _08656_ (.A(net517),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__mux4_1 _08657_ (.A0(\dpath.RF.R[16][12] ),
    .A1(\dpath.RF.R[17][12] ),
    .A2(\dpath.RF.R[18][12] ),
    .A3(\dpath.RF.R[19][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02863_));
 sky130_fd_sc_hd__nor2_1 _08658_ (.A(net533),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__mux4_1 _08659_ (.A0(\dpath.RF.R[20][12] ),
    .A1(\dpath.RF.R[21][12] ),
    .A2(\dpath.RF.R[22][12] ),
    .A3(\dpath.RF.R[23][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02865_));
 sky130_fd_sc_hd__nor2_1 _08660_ (.A(net509),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__mux4_1 _08661_ (.A0(\dpath.RF.R[28][12] ),
    .A1(\dpath.RF.R[29][12] ),
    .A2(\dpath.RF.R[30][12] ),
    .A3(\dpath.RF.R[31][12] ),
    .S0(net561),
    .S1(net542),
    .X(_02867_));
 sky130_fd_sc_hd__nor2_1 _08662_ (.A(net509),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__mux4_1 _08663_ (.A0(\dpath.RF.R[24][12] ),
    .A1(\dpath.RF.R[25][12] ),
    .A2(\dpath.RF.R[26][12] ),
    .A3(\dpath.RF.R[27][12] ),
    .S0(net560),
    .S1(net541),
    .X(_02869_));
 sky130_fd_sc_hd__o21ai_1 _08664_ (.A1(net530),
    .A2(_02869_),
    .B1(net522),
    .Y(_02870_));
 sky130_fd_sc_hd__o32a_1 _08665_ (.A1(net522),
    .A2(_02864_),
    .A3(_02866_),
    .B1(_02868_),
    .B2(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__a221o_1 _08666_ (.A1(_02857_),
    .A2(_02862_),
    .B1(_02871_),
    .B2(net517),
    .C1(net482),
    .X(_02872_));
 sky130_fd_sc_hd__nor2_1 _08667_ (.A(net372),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__mux2_2 _08668_ (.A0(net3638),
    .A1(net4),
    .S(net479),
    .X(_02874_));
 sky130_fd_sc_hd__a221o_1 _08669_ (.A1(net694),
    .A2(net370),
    .B1(net368),
    .B2(_02874_),
    .C1(_02873_),
    .X(_02875_));
 sky130_fd_sc_hd__nand2_1 _08670_ (.A(net632),
    .B(net757),
    .Y(_02876_));
 sky130_fd_sc_hd__a22oi_2 _08671_ (.A1(net636),
    .A2(net754),
    .B1(net751),
    .B2(net642),
    .Y(_02877_));
 sky130_fd_sc_hd__and4_1 _08672_ (.A(net642),
    .B(net637),
    .C(net754),
    .D(net751),
    .X(_02878_));
 sky130_fd_sc_hd__nor2_1 _08673_ (.A(_02877_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__xnor2_1 _08674_ (.A(_02876_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__a22o_1 _08675_ (.A1(net646),
    .A2(net748),
    .B1(net744),
    .B2(net651),
    .X(_02881_));
 sky130_fd_sc_hd__and4_1 _08676_ (.A(net650),
    .B(net647),
    .C(net748),
    .D(net744),
    .X(_02882_));
 sky130_fd_sc_hd__nand4_1 _08677_ (.A(net651),
    .B(net646),
    .C(net748),
    .D(net744),
    .Y(_02883_));
 sky130_fd_sc_hd__and3_1 _08678_ (.A(_02880_),
    .B(_02881_),
    .C(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__a21oi_1 _08679_ (.A1(_02881_),
    .A2(_02883_),
    .B1(_02880_),
    .Y(_02885_));
 sky130_fd_sc_hd__or2_1 _08680_ (.A(_02884_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__o21ba_1 _08681_ (.A1(_02789_),
    .A2(_02797_),
    .B1_N(_02796_),
    .X(_02887_));
 sky130_fd_sc_hd__nand2_1 _08682_ (.A(net785),
    .B(net608),
    .Y(_02888_));
 sky130_fd_sc_hd__and2_1 _08683_ (.A(net781),
    .B(net611),
    .X(_02889_));
 sky130_fd_sc_hd__a22o_1 _08684_ (.A1(net774),
    .A2(net617),
    .B1(net613),
    .B2(net779),
    .X(_02890_));
 sky130_fd_sc_hd__nand4_2 _08685_ (.A(net779),
    .B(net774),
    .C(net617),
    .D(net613),
    .Y(_02891_));
 sky130_fd_sc_hd__nand3_1 _08686_ (.A(_02889_),
    .B(_02890_),
    .C(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__a21o_1 _08687_ (.A1(_02890_),
    .A2(_02891_),
    .B1(_02889_),
    .X(_02893_));
 sky130_fd_sc_hd__a21bo_1 _08688_ (.A1(_02790_),
    .A2(_02791_),
    .B1_N(_02792_),
    .X(_02894_));
 sky130_fd_sc_hd__and3_1 _08689_ (.A(_02892_),
    .B(_02893_),
    .C(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__a21oi_1 _08690_ (.A1(_02892_),
    .A2(_02893_),
    .B1(_02894_),
    .Y(_02896_));
 sky130_fd_sc_hd__nor2_1 _08691_ (.A(_02895_),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__xnor2_1 _08692_ (.A(_02888_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2b_1 _08693_ (.A_N(_02887_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__xnor2_1 _08694_ (.A(_02887_),
    .B(_02898_),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(net788),
    .B(net606),
    .Y(_02901_));
 sky130_fd_sc_hd__nand3_1 _08696_ (.A(net788),
    .B(net606),
    .C(_02900_),
    .Y(_02902_));
 sky130_fd_sc_hd__xnor2_1 _08697_ (.A(_02900_),
    .B(_02901_),
    .Y(_02903_));
 sky130_fd_sc_hd__a32o_1 _08698_ (.A1(_02808_),
    .A2(_02811_),
    .A3(_02812_),
    .B1(_02814_),
    .B2(_02807_),
    .X(_02904_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(_02810_),
    .B(_02811_),
    .Y(_02905_));
 sky130_fd_sc_hd__a32o_1 _08700_ (.A1(net636),
    .A2(net757),
    .A3(_02780_),
    .B1(_02781_),
    .B2(net754),
    .X(_02906_));
 sky130_fd_sc_hd__a22o_1 _08701_ (.A1(net627),
    .A2(net765),
    .B1(net762),
    .B2(net628),
    .X(_02907_));
 sky130_fd_sc_hd__nand4_2 _08702_ (.A(net628),
    .B(net624),
    .C(net765),
    .D(net762),
    .Y(_02908_));
 sky130_fd_sc_hd__nand4_2 _08703_ (.A(net770),
    .B(net620),
    .C(_02907_),
    .D(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a22o_1 _08704_ (.A1(net770),
    .A2(net620),
    .B1(_02907_),
    .B2(_02908_),
    .X(_02910_));
 sky130_fd_sc_hd__nand3_1 _08705_ (.A(_02906_),
    .B(_02909_),
    .C(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21o_1 _08706_ (.A1(_02909_),
    .A2(_02910_),
    .B1(_02906_),
    .X(_02912_));
 sky130_fd_sc_hd__nand3_1 _08707_ (.A(_02905_),
    .B(_02911_),
    .C(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__a21o_1 _08708_ (.A1(_02911_),
    .A2(_02912_),
    .B1(_02905_),
    .X(_02914_));
 sky130_fd_sc_hd__nand3_1 _08709_ (.A(_02784_),
    .B(_02913_),
    .C(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__inv_2 _08710_ (.A(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__a21o_1 _08711_ (.A1(_02913_),
    .A2(_02914_),
    .B1(_02784_),
    .X(_02917_));
 sky130_fd_sc_hd__and3_2 _08712_ (.A(_02904_),
    .B(_02915_),
    .C(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__a21oi_1 _08713_ (.A1(_02915_),
    .A2(_02917_),
    .B1(_02904_),
    .Y(_02919_));
 sky130_fd_sc_hd__or3_4 _08714_ (.A(_02816_),
    .B(_02918_),
    .C(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__o21ai_2 _08715_ (.A1(_02918_),
    .A2(_02919_),
    .B1(_02816_),
    .Y(_02921_));
 sky130_fd_sc_hd__and3_1 _08716_ (.A(_02903_),
    .B(_02920_),
    .C(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__nand3_2 _08717_ (.A(_02903_),
    .B(_02920_),
    .C(_02921_),
    .Y(_02923_));
 sky130_fd_sc_hd__a21oi_1 _08718_ (.A1(_02920_),
    .A2(_02921_),
    .B1(_02903_),
    .Y(_02924_));
 sky130_fd_sc_hd__a211o_2 _08719_ (.A1(_02818_),
    .A2(_02820_),
    .B1(_02922_),
    .C1(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__o211ai_2 _08720_ (.A1(_02922_),
    .A2(_02924_),
    .B1(_02818_),
    .C1(_02820_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand3b_2 _08721_ (.A_N(_02886_),
    .B(_02925_),
    .C(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__a21bo_1 _08722_ (.A1(_02925_),
    .A2(_02926_),
    .B1_N(_02886_),
    .X(_02928_));
 sky130_fd_sc_hd__o211a_1 _08723_ (.A1(_02822_),
    .A2(_02824_),
    .B1(_02927_),
    .C1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__a211oi_2 _08724_ (.A1(_02927_),
    .A2(_02928_),
    .B1(_02822_),
    .C1(_02824_),
    .Y(_02930_));
 sky130_fd_sc_hd__or3b_4 _08725_ (.A(_02929_),
    .B(_02930_),
    .C_N(_02826_),
    .X(_02931_));
 sky130_fd_sc_hd__o21bai_2 _08726_ (.A1(_02929_),
    .A2(_02930_),
    .B1_N(_02826_),
    .Y(_02932_));
 sky130_fd_sc_hd__o211ai_4 _08727_ (.A1(_02800_),
    .A2(_02803_),
    .B1(_02931_),
    .C1(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__a211o_1 _08728_ (.A1(_02931_),
    .A2(_02932_),
    .B1(_02800_),
    .C1(_02803_),
    .X(_02934_));
 sky130_fd_sc_hd__o211ai_2 _08729_ (.A1(_02828_),
    .A2(_02830_),
    .B1(_02933_),
    .C1(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__a211o_1 _08730_ (.A1(_02933_),
    .A2(_02934_),
    .B1(_02828_),
    .C1(_02830_),
    .X(_02936_));
 sky130_fd_sc_hd__and2_1 _08731_ (.A(_02935_),
    .B(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__o21a_1 _08732_ (.A1(_02778_),
    .A2(_02834_),
    .B1(_02833_),
    .X(_02938_));
 sky130_fd_sc_hd__o311ai_4 _08733_ (.A1(_02728_),
    .A2(_02732_),
    .A3(_02834_),
    .B1(_02937_),
    .C1(_02833_),
    .Y(_02939_));
 sky130_fd_sc_hd__or2_1 _08734_ (.A(_02937_),
    .B(_02938_),
    .X(_02940_));
 sky130_fd_sc_hd__and3_1 _08735_ (.A(_02239_),
    .B(_02939_),
    .C(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__a21o_1 _08736_ (.A1(_01885_),
    .A2(_02777_),
    .B1(_01878_),
    .X(_02942_));
 sky130_fd_sc_hd__a31oi_1 _08737_ (.A1(_01878_),
    .A2(_01885_),
    .A3(_02777_),
    .B1(net468),
    .Y(_02943_));
 sky130_fd_sc_hd__a221o_4 _08738_ (.A1(net3346),
    .A2(net485),
    .B1(_02942_),
    .B2(_02943_),
    .C1(_02941_),
    .X(_02944_));
 sky130_fd_sc_hd__a21oi_4 _08739_ (.A1(net392),
    .A2(_02944_),
    .B1(_02875_),
    .Y(_02945_));
 sky130_fd_sc_hd__and2b_4 _08740_ (.A_N(_01836_),
    .B(net577),
    .X(_02946_));
 sky130_fd_sc_hd__and2_1 _08741_ (.A(net3264),
    .B(_01836_),
    .X(_02947_));
 sky130_fd_sc_hd__o21a_1 _08742_ (.A1(_02946_),
    .A2(_02947_),
    .B1(net3301),
    .X(_02948_));
 sky130_fd_sc_hd__or3_1 _08743_ (.A(net3301),
    .B(_02946_),
    .C(_02947_),
    .X(_02949_));
 sky130_fd_sc_hd__and2b_1 _08744_ (.A_N(_02948_),
    .B(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__a21o_1 _08745_ (.A1(_02847_),
    .A2(_02848_),
    .B1(_02846_),
    .X(_02951_));
 sky130_fd_sc_hd__xnor2_1 _08746_ (.A(_02950_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__o2bb2a_1 _08747_ (.A1_N(\dpath.btarg_DX.q[12] ),
    .A2_N(net403),
    .B1(net365),
    .B2(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__o211a_1 _08748_ (.A1(net373),
    .A2(_02945_),
    .B1(_02953_),
    .C1(_01958_),
    .X(_02954_));
 sky130_fd_sc_hd__a21oi_1 _08749_ (.A1(net361),
    .A2(_02853_),
    .B1(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__or2_1 _08750_ (.A(net3579),
    .B(net441),
    .X(_02956_));
 sky130_fd_sc_hd__o211a_1 _08751_ (.A1(net449),
    .A2(_02955_),
    .B1(_02956_),
    .C1(net845),
    .X(_00648_));
 sky130_fd_sc_hd__mux4_1 _08752_ (.A0(\dpath.RF.R[0][13] ),
    .A1(\dpath.RF.R[1][13] ),
    .A2(\dpath.RF.R[2][13] ),
    .A3(\dpath.RF.R[3][13] ),
    .S0(net559),
    .S1(net540),
    .X(_02957_));
 sky130_fd_sc_hd__mux4_1 _08753_ (.A0(\dpath.RF.R[4][13] ),
    .A1(\dpath.RF.R[5][13] ),
    .A2(\dpath.RF.R[6][13] ),
    .A3(\dpath.RF.R[7][13] ),
    .S0(net559),
    .S1(net540),
    .X(_02958_));
 sky130_fd_sc_hd__o21a_1 _08754_ (.A1(net509),
    .A2(_02958_),
    .B1(net506),
    .X(_02959_));
 sky130_fd_sc_hd__o21ai_1 _08755_ (.A1(net530),
    .A2(_02957_),
    .B1(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__mux4_1 _08756_ (.A0(\dpath.RF.R[12][13] ),
    .A1(\dpath.RF.R[13][13] ),
    .A2(\dpath.RF.R[14][13] ),
    .A3(\dpath.RF.R[15][13] ),
    .S0(net559),
    .S1(net540),
    .X(_02961_));
 sky130_fd_sc_hd__mux4_1 _08757_ (.A0(\dpath.RF.R[8][13] ),
    .A1(\dpath.RF.R[9][13] ),
    .A2(\dpath.RF.R[10][13] ),
    .A3(\dpath.RF.R[11][13] ),
    .S0(net561),
    .S1(net542),
    .X(_02962_));
 sky130_fd_sc_hd__or2_1 _08758_ (.A(net530),
    .B(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__o211a_1 _08759_ (.A1(net509),
    .A2(_02961_),
    .B1(_02963_),
    .C1(net522),
    .X(_02964_));
 sky130_fd_sc_hd__nor2_1 _08760_ (.A(net517),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__mux4_1 _08761_ (.A0(\dpath.RF.R[16][13] ),
    .A1(\dpath.RF.R[17][13] ),
    .A2(\dpath.RF.R[18][13] ),
    .A3(\dpath.RF.R[19][13] ),
    .S0(net561),
    .S1(net542),
    .X(_02966_));
 sky130_fd_sc_hd__nor2_1 _08762_ (.A(net530),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__mux4_1 _08763_ (.A0(\dpath.RF.R[20][13] ),
    .A1(\dpath.RF.R[21][13] ),
    .A2(\dpath.RF.R[22][13] ),
    .A3(\dpath.RF.R[23][13] ),
    .S0(net561),
    .S1(net542),
    .X(_02968_));
 sky130_fd_sc_hd__nor2_1 _08764_ (.A(net509),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__mux4_1 _08765_ (.A0(\dpath.RF.R[28][13] ),
    .A1(\dpath.RF.R[29][13] ),
    .A2(\dpath.RF.R[30][13] ),
    .A3(\dpath.RF.R[31][13] ),
    .S0(net559),
    .S1(net540),
    .X(_02970_));
 sky130_fd_sc_hd__nor2_1 _08766_ (.A(net509),
    .B(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__mux4_1 _08767_ (.A0(\dpath.RF.R[24][13] ),
    .A1(\dpath.RF.R[25][13] ),
    .A2(\dpath.RF.R[26][13] ),
    .A3(\dpath.RF.R[27][13] ),
    .S0(net559),
    .S1(net540),
    .X(_02972_));
 sky130_fd_sc_hd__o21ai_1 _08768_ (.A1(net530),
    .A2(_02972_),
    .B1(net522),
    .Y(_02973_));
 sky130_fd_sc_hd__o32a_1 _08769_ (.A1(net522),
    .A2(_02967_),
    .A3(_02969_),
    .B1(_02971_),
    .B2(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__a221o_1 _08770_ (.A1(_02960_),
    .A2(_02965_),
    .B1(_02974_),
    .B2(net517),
    .C1(net482),
    .X(_02975_));
 sky130_fd_sc_hd__nor2_1 _08771_ (.A(net372),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__mux2_1 _08772_ (.A0(net3621),
    .A1(net5),
    .S(net479),
    .X(_02977_));
 sky130_fd_sc_hd__a221o_1 _08773_ (.A1(net3586),
    .A2(net370),
    .B1(net368),
    .B2(_02977_),
    .C1(_02976_),
    .X(_02978_));
 sky130_fd_sc_hd__nand2_1 _08774_ (.A(net629),
    .B(net757),
    .Y(_02979_));
 sky130_fd_sc_hd__a22o_1 _08775_ (.A1(net632),
    .A2(net754),
    .B1(net751),
    .B2(net636),
    .X(_02980_));
 sky130_fd_sc_hd__and3_1 _08776_ (.A(net636),
    .B(net632),
    .C(net751),
    .X(_02981_));
 sky130_fd_sc_hd__a21bo_1 _08777_ (.A1(\dpath.alu.adder.in1[9] ),
    .A2(_02981_),
    .B1_N(_02980_),
    .X(_02982_));
 sky130_fd_sc_hd__xor2_2 _08778_ (.A(_02979_),
    .B(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__a22o_1 _08779_ (.A1(net647),
    .A2(net744),
    .B1(net740),
    .B2(net650),
    .X(_02984_));
 sky130_fd_sc_hd__and4_1 _08780_ (.A(net650),
    .B(net647),
    .C(net744),
    .D(net740),
    .X(_02985_));
 sky130_fd_sc_hd__nand4_1 _08781_ (.A(net650),
    .B(net647),
    .C(net744),
    .D(net740),
    .Y(_02986_));
 sky130_fd_sc_hd__and4_1 _08782_ (.A(net642),
    .B(net748),
    .C(_02984_),
    .D(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__nand4_1 _08783_ (.A(net642),
    .B(net748),
    .C(_02984_),
    .D(_02986_),
    .Y(_02988_));
 sky130_fd_sc_hd__a22o_1 _08784_ (.A1(net642),
    .A2(net748),
    .B1(_02984_),
    .B2(_02986_),
    .X(_02989_));
 sky130_fd_sc_hd__and3_1 _08785_ (.A(_02882_),
    .B(_02988_),
    .C(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__a21o_1 _08786_ (.A1(_02988_),
    .A2(_02989_),
    .B1(_02882_),
    .X(_02991_));
 sky130_fd_sc_hd__and2b_1 _08787_ (.A_N(_02990_),
    .B(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__xnor2_2 _08788_ (.A(_02983_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__o21ba_1 _08789_ (.A1(_02888_),
    .A2(_02896_),
    .B1_N(_02895_),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_1 _08790_ (.A(net785),
    .B(net606),
    .Y(_02995_));
 sky130_fd_sc_hd__and2_1 _08791_ (.A(net781),
    .B(net608),
    .X(_02996_));
 sky130_fd_sc_hd__a22o_1 _08792_ (.A1(net774),
    .A2(net613),
    .B1(net612),
    .B2(net779),
    .X(_02997_));
 sky130_fd_sc_hd__nand4_1 _08793_ (.A(net779),
    .B(net774),
    .C(net613),
    .D(net612),
    .Y(_02998_));
 sky130_fd_sc_hd__nand3_1 _08794_ (.A(_02996_),
    .B(_02997_),
    .C(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21o_1 _08795_ (.A1(_02997_),
    .A2(_02998_),
    .B1(_02996_),
    .X(_03000_));
 sky130_fd_sc_hd__a21bo_1 _08796_ (.A1(_02889_),
    .A2(_02890_),
    .B1_N(_02891_),
    .X(_03001_));
 sky130_fd_sc_hd__and3_1 _08797_ (.A(_02999_),
    .B(_03000_),
    .C(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__a21oi_1 _08798_ (.A1(_02999_),
    .A2(_03000_),
    .B1(_03001_),
    .Y(_03003_));
 sky130_fd_sc_hd__nor2_1 _08799_ (.A(_03002_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__xnor2_2 _08800_ (.A(_02995_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__and2b_1 _08801_ (.A_N(_02994_),
    .B(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__xnor2_2 _08802_ (.A(_02994_),
    .B(_03005_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _08803_ (.A(net788),
    .B(net603),
    .Y(_03008_));
 sky130_fd_sc_hd__xnor2_2 _08804_ (.A(_03007_),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_02911_),
    .B(_02913_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _08806_ (.A(_02908_),
    .B(_02909_),
    .Y(_03011_));
 sky130_fd_sc_hd__o21bai_2 _08807_ (.A1(_02876_),
    .A2(_02877_),
    .B1_N(_02878_),
    .Y(_03012_));
 sky130_fd_sc_hd__a22o_1 _08808_ (.A1(net765),
    .A2(net620),
    .B1(net762),
    .B2(net625),
    .X(_03013_));
 sky130_fd_sc_hd__nand4_2 _08809_ (.A(net625),
    .B(net765),
    .C(net621),
    .D(net762),
    .Y(_03014_));
 sky130_fd_sc_hd__nand4_2 _08810_ (.A(net770),
    .B(net616),
    .C(_03013_),
    .D(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__a22o_1 _08811_ (.A1(net770),
    .A2(net616),
    .B1(_03013_),
    .B2(_03014_),
    .X(_03016_));
 sky130_fd_sc_hd__nand3_2 _08812_ (.A(_03012_),
    .B(_03015_),
    .C(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__a21o_1 _08813_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03012_),
    .X(_03018_));
 sky130_fd_sc_hd__nand3_2 _08814_ (.A(_03011_),
    .B(_03017_),
    .C(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__a21o_1 _08815_ (.A1(_03017_),
    .A2(_03018_),
    .B1(_03011_),
    .X(_03020_));
 sky130_fd_sc_hd__nand3_2 _08816_ (.A(_02884_),
    .B(_03019_),
    .C(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__inv_2 _08817_ (.A(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__a21o_1 _08818_ (.A1(_03019_),
    .A2(_03020_),
    .B1(_02884_),
    .X(_03023_));
 sky130_fd_sc_hd__and3_1 _08819_ (.A(_03010_),
    .B(_03021_),
    .C(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__nand3_2 _08820_ (.A(_03010_),
    .B(_03021_),
    .C(_03023_),
    .Y(_03025_));
 sky130_fd_sc_hd__a21o_1 _08821_ (.A1(_03021_),
    .A2(_03023_),
    .B1(_03010_),
    .X(_03026_));
 sky130_fd_sc_hd__o211ai_4 _08822_ (.A1(_02916_),
    .A2(_02918_),
    .B1(_03025_),
    .C1(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__a211o_1 _08823_ (.A1(_03025_),
    .A2(_03026_),
    .B1(_02916_),
    .C1(_02918_),
    .X(_03028_));
 sky130_fd_sc_hd__and3_1 _08824_ (.A(_03009_),
    .B(_03027_),
    .C(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__nand3_2 _08825_ (.A(_03009_),
    .B(_03027_),
    .C(_03028_),
    .Y(_03030_));
 sky130_fd_sc_hd__a21oi_2 _08826_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_03009_),
    .Y(_03031_));
 sky130_fd_sc_hd__a211oi_4 _08827_ (.A1(_02920_),
    .A2(_02923_),
    .B1(_03029_),
    .C1(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__o211a_1 _08828_ (.A1(_03029_),
    .A2(_03031_),
    .B1(_02920_),
    .C1(_02923_),
    .X(_03033_));
 sky130_fd_sc_hd__nor3_2 _08829_ (.A(_02993_),
    .B(_03032_),
    .C(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__o21a_1 _08830_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_02993_),
    .X(_03035_));
 sky130_fd_sc_hd__a211oi_2 _08831_ (.A1(_02925_),
    .A2(_02927_),
    .B1(_03034_),
    .C1(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__o211a_1 _08832_ (.A1(_03034_),
    .A2(_03035_),
    .B1(_02925_),
    .C1(_02927_),
    .X(_03037_));
 sky130_fd_sc_hd__nor3b_1 _08833_ (.A(_03036_),
    .B(_03037_),
    .C_N(_02929_),
    .Y(_03038_));
 sky130_fd_sc_hd__o21ba_1 _08834_ (.A1(_03036_),
    .A2(_03037_),
    .B1_N(_02929_),
    .X(_03039_));
 sky130_fd_sc_hd__a211oi_2 _08835_ (.A1(_02899_),
    .A2(_02902_),
    .B1(_03038_),
    .C1(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__o211a_1 _08836_ (.A1(_03038_),
    .A2(_03039_),
    .B1(_02899_),
    .C1(_02902_),
    .X(_03041_));
 sky130_fd_sc_hd__a211oi_1 _08837_ (.A1(_02931_),
    .A2(_02933_),
    .B1(_03040_),
    .C1(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__a211o_1 _08838_ (.A1(_02931_),
    .A2(_02933_),
    .B1(_03040_),
    .C1(_03041_),
    .X(_03043_));
 sky130_fd_sc_hd__o211a_1 _08839_ (.A1(_03040_),
    .A2(_03041_),
    .B1(_02931_),
    .C1(_02933_),
    .X(_03044_));
 sky130_fd_sc_hd__nor2_1 _08840_ (.A(_03042_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_02935_),
    .B(_02939_),
    .Y(_03046_));
 sky130_fd_sc_hd__xor2_1 _08842_ (.A(_03045_),
    .B(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__or2_1 _08843_ (.A(net3688),
    .B(net484),
    .X(_03048_));
 sky130_fd_sc_hd__o211a_1 _08844_ (.A1(net485),
    .A2(_03047_),
    .B1(_03048_),
    .C1(net468),
    .X(_03049_));
 sky130_fd_sc_hd__a21bo_1 _08845_ (.A1(_01876_),
    .A2(_02942_),
    .B1_N(_01850_),
    .X(_03050_));
 sky130_fd_sc_hd__nand3b_1 _08846_ (.A_N(_01850_),
    .B(_01876_),
    .C(_02942_),
    .Y(_03051_));
 sky130_fd_sc_hd__a31o_4 _08847_ (.A1(net467),
    .A2(_03050_),
    .A3(_03051_),
    .B1(_03049_),
    .X(_03052_));
 sky130_fd_sc_hd__a21o_4 _08848_ (.A1(net392),
    .A2(_03052_),
    .B1(_02978_),
    .X(_03053_));
 sky130_fd_sc_hd__and2_1 _08849_ (.A(net3282),
    .B(_01836_),
    .X(_03054_));
 sky130_fd_sc_hd__o21a_1 _08850_ (.A1(_02946_),
    .A2(_03054_),
    .B1(net3295),
    .X(_03055_));
 sky130_fd_sc_hd__or3_1 _08851_ (.A(net3295),
    .B(_02946_),
    .C(_03054_),
    .X(_03056_));
 sky130_fd_sc_hd__and2b_1 _08852_ (.A_N(_03055_),
    .B(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__a21o_1 _08853_ (.A1(_02949_),
    .A2(_02951_),
    .B1(_02948_),
    .X(_03058_));
 sky130_fd_sc_hd__xnor2_1 _08854_ (.A(_03057_),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__a21oi_1 _08855_ (.A1(net231),
    .A2(_02751_),
    .B1(net3539),
    .Y(_03060_));
 sky130_fd_sc_hd__and3_1 _08856_ (.A(net3539),
    .B(net231),
    .C(_02751_),
    .X(_03061_));
 sky130_fd_sc_hd__or3_1 _08857_ (.A(_01958_),
    .B(_03060_),
    .C(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__a21oi_1 _08858_ (.A1(\dpath.btarg_DX.q[13] ),
    .A2(net403),
    .B1(net449),
    .Y(_03063_));
 sky130_fd_sc_hd__o211a_1 _08859_ (.A1(net365),
    .A2(_03059_),
    .B1(_03062_),
    .C1(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__a21bo_1 _08860_ (.A1(_02027_),
    .A2(_03053_),
    .B1_N(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__o211a_1 _08861_ (.A1(net3539),
    .A2(net441),
    .B1(_03065_),
    .C1(net845),
    .X(_00649_));
 sky130_fd_sc_hd__xnor2_1 _08862_ (.A(net3555),
    .B(_03061_),
    .Y(_03066_));
 sky130_fd_sc_hd__mux4_1 _08863_ (.A0(\dpath.RF.R[0][14] ),
    .A1(\dpath.RF.R[1][14] ),
    .A2(\dpath.RF.R[2][14] ),
    .A3(\dpath.RF.R[3][14] ),
    .S0(net560),
    .S1(net541),
    .X(_03067_));
 sky130_fd_sc_hd__mux4_1 _08864_ (.A0(\dpath.RF.R[4][14] ),
    .A1(\dpath.RF.R[5][14] ),
    .A2(\dpath.RF.R[6][14] ),
    .A3(\dpath.RF.R[7][14] ),
    .S0(net560),
    .S1(net541),
    .X(_03068_));
 sky130_fd_sc_hd__o21a_1 _08865_ (.A1(net509),
    .A2(_03068_),
    .B1(net506),
    .X(_03069_));
 sky130_fd_sc_hd__o21ai_1 _08866_ (.A1(net530),
    .A2(_03067_),
    .B1(_03069_),
    .Y(_03070_));
 sky130_fd_sc_hd__mux4_1 _08867_ (.A0(\dpath.RF.R[12][14] ),
    .A1(\dpath.RF.R[13][14] ),
    .A2(\dpath.RF.R[14][14] ),
    .A3(\dpath.RF.R[15][14] ),
    .S0(net567),
    .S1(net548),
    .X(_03071_));
 sky130_fd_sc_hd__mux4_1 _08868_ (.A0(\dpath.RF.R[8][14] ),
    .A1(\dpath.RF.R[9][14] ),
    .A2(\dpath.RF.R[10][14] ),
    .A3(\dpath.RF.R[11][14] ),
    .S0(net560),
    .S1(net541),
    .X(_03072_));
 sky130_fd_sc_hd__or2_1 _08869_ (.A(net533),
    .B(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__o211a_1 _08870_ (.A1(net510),
    .A2(_03071_),
    .B1(_03073_),
    .C1(net522),
    .X(_03074_));
 sky130_fd_sc_hd__nor2_1 _08871_ (.A(_00009_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__mux4_1 _08872_ (.A0(\dpath.RF.R[16][14] ),
    .A1(\dpath.RF.R[17][14] ),
    .A2(\dpath.RF.R[18][14] ),
    .A3(\dpath.RF.R[19][14] ),
    .S0(net571),
    .S1(net552),
    .X(_03076_));
 sky130_fd_sc_hd__nor2_1 _08873_ (.A(net532),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__mux4_1 _08874_ (.A0(\dpath.RF.R[20][14] ),
    .A1(\dpath.RF.R[21][14] ),
    .A2(\dpath.RF.R[22][14] ),
    .A3(\dpath.RF.R[23][14] ),
    .S0(net565),
    .S1(net544),
    .X(_03078_));
 sky130_fd_sc_hd__nor2_1 _08875_ (.A(net512),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__mux4_1 _08876_ (.A0(\dpath.RF.R[28][14] ),
    .A1(\dpath.RF.R[29][14] ),
    .A2(\dpath.RF.R[30][14] ),
    .A3(\dpath.RF.R[31][14] ),
    .S0(net571),
    .S1(net552),
    .X(_03080_));
 sky130_fd_sc_hd__nor2_1 _08877_ (.A(net512),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__mux4_1 _08878_ (.A0(\dpath.RF.R[24][14] ),
    .A1(\dpath.RF.R[25][14] ),
    .A2(\dpath.RF.R[26][14] ),
    .A3(\dpath.RF.R[27][14] ),
    .S0(net565),
    .S1(net544),
    .X(_03082_));
 sky130_fd_sc_hd__o21ai_1 _08879_ (.A1(net532),
    .A2(_03082_),
    .B1(net524),
    .Y(_03083_));
 sky130_fd_sc_hd__o32a_1 _08880_ (.A1(net524),
    .A2(_03077_),
    .A3(_03079_),
    .B1(_03081_),
    .B2(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__a221o_1 _08881_ (.A1(_03070_),
    .A2(_03075_),
    .B1(_03084_),
    .B2(net518),
    .C1(net482),
    .X(_03085_));
 sky130_fd_sc_hd__nor2_1 _08882_ (.A(net371),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__mux2_2 _08883_ (.A0(net3639),
    .A1(net6),
    .S(net479),
    .X(_03087_));
 sky130_fd_sc_hd__a221o_1 _08884_ (.A1(net691),
    .A2(net369),
    .B1(net367),
    .B2(_03087_),
    .C1(_03086_),
    .X(_03088_));
 sky130_fd_sc_hd__a31o_1 _08885_ (.A1(net788),
    .A2(net603),
    .A3(_03007_),
    .B1(_03006_),
    .X(_03089_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(net625),
    .B(net757),
    .Y(_03090_));
 sky130_fd_sc_hd__a22o_1 _08887_ (.A1(net629),
    .A2(net754),
    .B1(net751),
    .B2(net633),
    .X(_03091_));
 sky130_fd_sc_hd__and3_1 _08888_ (.A(net633),
    .B(net629),
    .C(net751),
    .X(_03092_));
 sky130_fd_sc_hd__a21bo_1 _08889_ (.A1(net754),
    .A2(_03092_),
    .B1_N(_03091_),
    .X(_03093_));
 sky130_fd_sc_hd__xor2_1 _08890_ (.A(_03090_),
    .B(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__a22o_1 _08891_ (.A1(net641),
    .A2(net744),
    .B1(net740),
    .B2(net646),
    .X(_03095_));
 sky130_fd_sc_hd__and4_1 _08892_ (.A(net647),
    .B(net641),
    .C(net744),
    .D(net740),
    .X(_03096_));
 sky130_fd_sc_hd__nand4_2 _08893_ (.A(net646),
    .B(net642),
    .C(net744),
    .D(net740),
    .Y(_03097_));
 sky130_fd_sc_hd__and4_1 _08894_ (.A(net637),
    .B(net748),
    .C(_03095_),
    .D(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__nand4_1 _08895_ (.A(net637),
    .B(net748),
    .C(_03095_),
    .D(_03097_),
    .Y(_03099_));
 sky130_fd_sc_hd__a22o_1 _08896_ (.A1(net637),
    .A2(net748),
    .B1(_03095_),
    .B2(_03097_),
    .X(_03100_));
 sky130_fd_sc_hd__o211a_1 _08897_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03099_),
    .C1(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__a211o_1 _08898_ (.A1(_03099_),
    .A2(_03100_),
    .B1(_02985_),
    .C1(_02987_),
    .X(_03102_));
 sky130_fd_sc_hd__and2b_1 _08899_ (.A_N(_03101_),
    .B(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__xor2_1 _08900_ (.A(_03094_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__nand3_1 _08901_ (.A(net650),
    .B(net736),
    .C(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__a21o_1 _08902_ (.A1(net650),
    .A2(net736),
    .B1(_03104_),
    .X(_03106_));
 sky130_fd_sc_hd__and2_1 _08903_ (.A(_03105_),
    .B(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__o21ba_1 _08904_ (.A1(_02995_),
    .A2(_03003_),
    .B1_N(_03002_),
    .X(_03108_));
 sky130_fd_sc_hd__nand2_1 _08905_ (.A(net785),
    .B(net603),
    .Y(_03109_));
 sky130_fd_sc_hd__and2_1 _08906_ (.A(net781),
    .B(net606),
    .X(_03110_));
 sky130_fd_sc_hd__a22o_1 _08907_ (.A1(net774),
    .A2(net612),
    .B1(net608),
    .B2(net779),
    .X(_03111_));
 sky130_fd_sc_hd__nand4_2 _08908_ (.A(net779),
    .B(net774),
    .C(net612),
    .D(net608),
    .Y(_03112_));
 sky130_fd_sc_hd__nand3_1 _08909_ (.A(_03110_),
    .B(_03111_),
    .C(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__a21o_1 _08910_ (.A1(_03111_),
    .A2(_03112_),
    .B1(_03110_),
    .X(_03114_));
 sky130_fd_sc_hd__a21bo_1 _08911_ (.A1(_02996_),
    .A2(_02997_),
    .B1_N(_02998_),
    .X(_03115_));
 sky130_fd_sc_hd__and3_1 _08912_ (.A(_03113_),
    .B(_03114_),
    .C(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__a21oi_1 _08913_ (.A1(_03113_),
    .A2(_03114_),
    .B1(_03115_),
    .Y(_03117_));
 sky130_fd_sc_hd__nor2_1 _08914_ (.A(_03116_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__xnor2_2 _08915_ (.A(_03109_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__and2b_1 _08916_ (.A_N(_03108_),
    .B(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__xnor2_2 _08917_ (.A(_03108_),
    .B(_03119_),
    .Y(_03121_));
 sky130_fd_sc_hd__nand2_1 _08918_ (.A(net788),
    .B(net600),
    .Y(_03122_));
 sky130_fd_sc_hd__and3_1 _08919_ (.A(net788),
    .B(net600),
    .C(_03121_),
    .X(_03123_));
 sky130_fd_sc_hd__xnor2_2 _08920_ (.A(_03121_),
    .B(_03122_),
    .Y(_03124_));
 sky130_fd_sc_hd__a21o_1 _08921_ (.A1(_02983_),
    .A2(_02991_),
    .B1(_02990_),
    .X(_03125_));
 sky130_fd_sc_hd__nand2_1 _08922_ (.A(_03014_),
    .B(_03015_),
    .Y(_03126_));
 sky130_fd_sc_hd__a32o_1 _08923_ (.A1(net629),
    .A2(net757),
    .A3(_02980_),
    .B1(_02981_),
    .B2(\dpath.alu.adder.in1[9] ),
    .X(_03127_));
 sky130_fd_sc_hd__a22o_1 _08924_ (.A1(net621),
    .A2(net763),
    .B1(net616),
    .B2(net765),
    .X(_03128_));
 sky130_fd_sc_hd__nand4_2 _08925_ (.A(net766),
    .B(net621),
    .C(net763),
    .D(net616),
    .Y(_03129_));
 sky130_fd_sc_hd__nand4_2 _08926_ (.A(net770),
    .B(net613),
    .C(_03128_),
    .D(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__a22o_1 _08927_ (.A1(net771),
    .A2(net613),
    .B1(_03128_),
    .B2(_03129_),
    .X(_03131_));
 sky130_fd_sc_hd__nand3_2 _08928_ (.A(_03127_),
    .B(_03130_),
    .C(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__a21o_1 _08929_ (.A1(_03130_),
    .A2(_03131_),
    .B1(_03127_),
    .X(_03133_));
 sky130_fd_sc_hd__nand3_2 _08930_ (.A(_03126_),
    .B(_03132_),
    .C(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__a21o_1 _08931_ (.A1(_03132_),
    .A2(_03133_),
    .B1(_03126_),
    .X(_03135_));
 sky130_fd_sc_hd__and3_2 _08932_ (.A(_03125_),
    .B(_03134_),
    .C(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__inv_2 _08933_ (.A(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__a21oi_2 _08934_ (.A1(_03134_),
    .A2(_03135_),
    .B1(_03125_),
    .Y(_03138_));
 sky130_fd_sc_hd__a211o_2 _08935_ (.A1(_03017_),
    .A2(_03019_),
    .B1(_03136_),
    .C1(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__o211ai_4 _08936_ (.A1(_03136_),
    .A2(_03138_),
    .B1(_03017_),
    .C1(_03019_),
    .Y(_03140_));
 sky130_fd_sc_hd__o211ai_4 _08937_ (.A1(_03022_),
    .A2(_03024_),
    .B1(_03139_),
    .C1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__a211o_1 _08938_ (.A1(_03139_),
    .A2(_03140_),
    .B1(_03022_),
    .C1(_03024_),
    .X(_03142_));
 sky130_fd_sc_hd__and3_1 _08939_ (.A(_03124_),
    .B(_03141_),
    .C(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__nand3_2 _08940_ (.A(_03124_),
    .B(_03141_),
    .C(_03142_),
    .Y(_03144_));
 sky130_fd_sc_hd__a21oi_2 _08941_ (.A1(_03141_),
    .A2(_03142_),
    .B1(_03124_),
    .Y(_03145_));
 sky130_fd_sc_hd__a211o_2 _08942_ (.A1(_03027_),
    .A2(_03030_),
    .B1(_03143_),
    .C1(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__o211ai_4 _08943_ (.A1(_03143_),
    .A2(_03145_),
    .B1(_03027_),
    .C1(_03030_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand3_4 _08944_ (.A(_03107_),
    .B(_03146_),
    .C(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__a21o_1 _08945_ (.A1(_03146_),
    .A2(_03147_),
    .B1(_03107_),
    .X(_03149_));
 sky130_fd_sc_hd__o211ai_4 _08946_ (.A1(_03032_),
    .A2(_03034_),
    .B1(_03148_),
    .C1(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__a211o_1 _08947_ (.A1(_03148_),
    .A2(_03149_),
    .B1(_03032_),
    .C1(_03034_),
    .X(_03151_));
 sky130_fd_sc_hd__nand3_2 _08948_ (.A(_03036_),
    .B(_03150_),
    .C(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__a21o_1 _08949_ (.A1(_03150_),
    .A2(_03151_),
    .B1(_03036_),
    .X(_03153_));
 sky130_fd_sc_hd__nand3_1 _08950_ (.A(_03089_),
    .B(_03152_),
    .C(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__a21o_1 _08951_ (.A1(_03152_),
    .A2(_03153_),
    .B1(_03089_),
    .X(_03155_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_03154_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__or2_1 _08953_ (.A(_03038_),
    .B(_03040_),
    .X(_03157_));
 sky130_fd_sc_hd__and3_1 _08954_ (.A(_03154_),
    .B(_03155_),
    .C(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__xnor2_2 _08955_ (.A(_03156_),
    .B(_03157_),
    .Y(_03159_));
 sky130_fd_sc_hd__o21ba_1 _08956_ (.A1(_03042_),
    .A2(_03046_),
    .B1_N(_03044_),
    .X(_03160_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__o211a_1 _08958_ (.A1(_03159_),
    .A2(_03160_),
    .B1(_03161_),
    .C1(_02239_),
    .X(_03162_));
 sky130_fd_sc_hd__a21o_1 _08959_ (.A1(_01848_),
    .A2(_03050_),
    .B1(_01897_),
    .X(_03163_));
 sky130_fd_sc_hd__a31o_1 _08960_ (.A1(_01848_),
    .A2(_01897_),
    .A3(_03050_),
    .B1(net468),
    .X(_03164_));
 sky130_fd_sc_hd__and2b_1 _08961_ (.A_N(_03164_),
    .B(_03163_),
    .X(_03165_));
 sky130_fd_sc_hd__a211o_4 _08962_ (.A1(net3504),
    .A2(net485),
    .B1(_03162_),
    .C1(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__a21oi_4 _08963_ (.A1(net391),
    .A2(_03166_),
    .B1(_03088_),
    .Y(_03167_));
 sky130_fd_sc_hd__and2_1 _08964_ (.A(net3342),
    .B(_02126_),
    .X(_03168_));
 sky130_fd_sc_hd__o21a_1 _08965_ (.A1(_02946_),
    .A2(_03168_),
    .B1(net3291),
    .X(_03169_));
 sky130_fd_sc_hd__or3_1 _08966_ (.A(net3291),
    .B(_02946_),
    .C(_03168_),
    .X(_03170_));
 sky130_fd_sc_hd__and2b_1 _08967_ (.A_N(_03169_),
    .B(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__a21o_1 _08968_ (.A1(_03056_),
    .A2(_03058_),
    .B1(_03055_),
    .X(_03172_));
 sky130_fd_sc_hd__xnor2_1 _08969_ (.A(_03171_),
    .B(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__o2bb2a_1 _08970_ (.A1_N(\dpath.btarg_DX.q[14] ),
    .A2_N(net403),
    .B1(net365),
    .B2(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__o211a_1 _08971_ (.A1(net373),
    .A2(_03167_),
    .B1(_03174_),
    .C1(_01958_),
    .X(_03175_));
 sky130_fd_sc_hd__a21oi_1 _08972_ (.A1(net361),
    .A2(_03066_),
    .B1(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__or2_1 _08973_ (.A(net3555),
    .B(net441),
    .X(_03177_));
 sky130_fd_sc_hd__o211a_1 _08974_ (.A1(net449),
    .A2(_03176_),
    .B1(_03177_),
    .C1(net845),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_1 _08975_ (.A0(\dpath.RF.R[0][15] ),
    .A1(\dpath.RF.R[1][15] ),
    .A2(\dpath.RF.R[2][15] ),
    .A3(\dpath.RF.R[3][15] ),
    .S0(net559),
    .S1(net540),
    .X(_03178_));
 sky130_fd_sc_hd__mux4_1 _08976_ (.A0(\dpath.RF.R[4][15] ),
    .A1(\dpath.RF.R[5][15] ),
    .A2(\dpath.RF.R[6][15] ),
    .A3(\dpath.RF.R[7][15] ),
    .S0(net559),
    .S1(net540),
    .X(_03179_));
 sky130_fd_sc_hd__o21a_1 _08977_ (.A1(net509),
    .A2(_03179_),
    .B1(net506),
    .X(_03180_));
 sky130_fd_sc_hd__o21ai_1 _08978_ (.A1(net530),
    .A2(_03178_),
    .B1(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__mux4_1 _08979_ (.A0(\dpath.RF.R[12][15] ),
    .A1(\dpath.RF.R[13][15] ),
    .A2(\dpath.RF.R[14][15] ),
    .A3(\dpath.RF.R[15][15] ),
    .S0(net566),
    .S1(net547),
    .X(_03182_));
 sky130_fd_sc_hd__mux4_1 _08980_ (.A0(\dpath.RF.R[8][15] ),
    .A1(\dpath.RF.R[9][15] ),
    .A2(\dpath.RF.R[10][15] ),
    .A3(\dpath.RF.R[11][15] ),
    .S0(net559),
    .S1(net540),
    .X(_03183_));
 sky130_fd_sc_hd__or2_1 _08981_ (.A(net530),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _08982_ (.A1(net509),
    .A2(_03182_),
    .B1(_03184_),
    .C1(net522),
    .X(_03185_));
 sky130_fd_sc_hd__nor2_1 _08983_ (.A(net518),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__mux4_1 _08984_ (.A0(\dpath.RF.R[16][15] ),
    .A1(\dpath.RF.R[17][15] ),
    .A2(\dpath.RF.R[18][15] ),
    .A3(\dpath.RF.R[19][15] ),
    .S0(net566),
    .S1(net547),
    .X(_03187_));
 sky130_fd_sc_hd__nor2_1 _08985_ (.A(net535),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__mux4_1 _08986_ (.A0(\dpath.RF.R[20][15] ),
    .A1(\dpath.RF.R[21][15] ),
    .A2(\dpath.RF.R[22][15] ),
    .A3(\dpath.RF.R[23][15] ),
    .S0(net559),
    .S1(net540),
    .X(_03189_));
 sky130_fd_sc_hd__nor2_1 _08987_ (.A(net509),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__mux4_1 _08988_ (.A0(\dpath.RF.R[28][15] ),
    .A1(\dpath.RF.R[29][15] ),
    .A2(\dpath.RF.R[30][15] ),
    .A3(\dpath.RF.R[31][15] ),
    .S0(net570),
    .S1(net551),
    .X(_03191_));
 sky130_fd_sc_hd__nor2_1 _08989_ (.A(net509),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__mux4_1 _08990_ (.A0(\dpath.RF.R[24][15] ),
    .A1(\dpath.RF.R[25][15] ),
    .A2(\dpath.RF.R[26][15] ),
    .A3(\dpath.RF.R[27][15] ),
    .S0(net559),
    .S1(net540),
    .X(_03193_));
 sky130_fd_sc_hd__o21ai_1 _08991_ (.A1(net530),
    .A2(_03193_),
    .B1(net522),
    .Y(_03194_));
 sky130_fd_sc_hd__o32a_1 _08992_ (.A1(net522),
    .A2(_03188_),
    .A3(_03190_),
    .B1(_03192_),
    .B2(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__a221o_1 _08993_ (.A1(_03181_),
    .A2(_03186_),
    .B1(_03195_),
    .B2(net518),
    .C1(net482),
    .X(_03196_));
 sky130_fd_sc_hd__nor2_1 _08994_ (.A(net371),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(net3634),
    .A1(net7),
    .S(net479),
    .X(_03198_));
 sky130_fd_sc_hd__a221o_1 _08996_ (.A1(net689),
    .A2(net369),
    .B1(net367),
    .B2(_03198_),
    .C1(_03197_),
    .X(_03199_));
 sky130_fd_sc_hd__nand2_2 _08997_ (.A(_03152_),
    .B(_03154_),
    .Y(_03200_));
 sky130_fd_sc_hd__a22o_1 _08998_ (.A1(net649),
    .A2(net736),
    .B1(net734),
    .B2(net653),
    .X(_03201_));
 sky130_fd_sc_hd__and3_1 _08999_ (.A(net652),
    .B(net649),
    .C(net734),
    .X(_03202_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(net736),
    .B(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(_03201_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nand2_1 _09002_ (.A(net621),
    .B(net758),
    .Y(_03205_));
 sky130_fd_sc_hd__a22o_1 _09003_ (.A1(net625),
    .A2(net755),
    .B1(net752),
    .B2(net629),
    .X(_03206_));
 sky130_fd_sc_hd__and3_1 _09004_ (.A(net629),
    .B(net625),
    .C(net752),
    .X(_03207_));
 sky130_fd_sc_hd__a21bo_1 _09005_ (.A1(net755),
    .A2(_03207_),
    .B1_N(_03206_),
    .X(_03208_));
 sky130_fd_sc_hd__xor2_1 _09006_ (.A(_03205_),
    .B(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__a22o_1 _09007_ (.A1(net637),
    .A2(net745),
    .B1(net740),
    .B2(net642),
    .X(_03210_));
 sky130_fd_sc_hd__and4_1 _09008_ (.A(net641),
    .B(net637),
    .C(net745),
    .D(net741),
    .X(_03211_));
 sky130_fd_sc_hd__nand4_1 _09009_ (.A(net642),
    .B(net637),
    .C(net744),
    .D(net740),
    .Y(_03212_));
 sky130_fd_sc_hd__and4_1 _09010_ (.A(net633),
    .B(net749),
    .C(_03210_),
    .D(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__nand4_1 _09011_ (.A(net633),
    .B(net749),
    .C(_03210_),
    .D(_03212_),
    .Y(_03214_));
 sky130_fd_sc_hd__a22o_1 _09012_ (.A1(net633),
    .A2(net749),
    .B1(_03210_),
    .B2(_03212_),
    .X(_03215_));
 sky130_fd_sc_hd__o211a_1 _09013_ (.A1(_03096_),
    .A2(_03098_),
    .B1(_03214_),
    .C1(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__a211o_1 _09014_ (.A1(_03214_),
    .A2(_03215_),
    .B1(_03096_),
    .C1(_03098_),
    .X(_03217_));
 sky130_fd_sc_hd__and2b_1 _09015_ (.A_N(_03216_),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__xnor2_1 _09016_ (.A(_03209_),
    .B(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__or2_1 _09017_ (.A(_03204_),
    .B(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__nand2_1 _09018_ (.A(_03204_),
    .B(_03219_),
    .Y(_03221_));
 sky130_fd_sc_hd__and2_1 _09019_ (.A(_03220_),
    .B(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__and2b_1 _09020_ (.A_N(_03105_),
    .B(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__xnor2_1 _09021_ (.A(_03105_),
    .B(_03222_),
    .Y(_03224_));
 sky130_fd_sc_hd__o21ba_1 _09022_ (.A1(_03109_),
    .A2(_03117_),
    .B1_N(_03116_),
    .X(_03225_));
 sky130_fd_sc_hd__nand2_1 _09023_ (.A(net785),
    .B(net600),
    .Y(_03226_));
 sky130_fd_sc_hd__and2_1 _09024_ (.A(net781),
    .B(net603),
    .X(_03227_));
 sky130_fd_sc_hd__a22o_1 _09025_ (.A1(net774),
    .A2(net608),
    .B1(net606),
    .B2(net779),
    .X(_03228_));
 sky130_fd_sc_hd__nand4_2 _09026_ (.A(net778),
    .B(net774),
    .C(net608),
    .D(net606),
    .Y(_03229_));
 sky130_fd_sc_hd__nand3_1 _09027_ (.A(_03227_),
    .B(_03228_),
    .C(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__a21o_1 _09028_ (.A1(_03228_),
    .A2(_03229_),
    .B1(_03227_),
    .X(_03231_));
 sky130_fd_sc_hd__a21bo_1 _09029_ (.A1(_03110_),
    .A2(_03111_),
    .B1_N(_03112_),
    .X(_03232_));
 sky130_fd_sc_hd__and3_1 _09030_ (.A(_03230_),
    .B(_03231_),
    .C(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__a21oi_1 _09031_ (.A1(_03230_),
    .A2(_03231_),
    .B1(_03232_),
    .Y(_03234_));
 sky130_fd_sc_hd__nor2_1 _09032_ (.A(_03233_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__xnor2_1 _09033_ (.A(_03226_),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__and2b_1 _09034_ (.A_N(_03225_),
    .B(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__xnor2_1 _09035_ (.A(_03225_),
    .B(_03236_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(net788),
    .B(net597),
    .Y(_03239_));
 sky130_fd_sc_hd__xnor2_1 _09037_ (.A(_03238_),
    .B(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__a21o_1 _09038_ (.A1(_03094_),
    .A2(_03102_),
    .B1(_03101_),
    .X(_03241_));
 sky130_fd_sc_hd__nand2_1 _09039_ (.A(_03129_),
    .B(_03130_),
    .Y(_03242_));
 sky130_fd_sc_hd__a32o_1 _09040_ (.A1(net625),
    .A2(net757),
    .A3(_03091_),
    .B1(_03092_),
    .B2(net754),
    .X(_03243_));
 sky130_fd_sc_hd__a22o_1 _09041_ (.A1(net761),
    .A2(net616),
    .B1(net615),
    .B2(net766),
    .X(_03244_));
 sky130_fd_sc_hd__nand4_2 _09042_ (.A(net766),
    .B(net761),
    .C(net616),
    .D(net615),
    .Y(_03245_));
 sky130_fd_sc_hd__nand4_2 _09043_ (.A(net769),
    .B(net611),
    .C(_03244_),
    .D(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__a22o_1 _09044_ (.A1(net769),
    .A2(net611),
    .B1(_03244_),
    .B2(_03245_),
    .X(_03247_));
 sky130_fd_sc_hd__nand3_4 _09045_ (.A(_03243_),
    .B(_03246_),
    .C(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__a21o_1 _09046_ (.A1(_03246_),
    .A2(_03247_),
    .B1(_03243_),
    .X(_03249_));
 sky130_fd_sc_hd__nand3_2 _09047_ (.A(_03242_),
    .B(_03248_),
    .C(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__a21o_1 _09048_ (.A1(_03248_),
    .A2(_03249_),
    .B1(_03242_),
    .X(_03251_));
 sky130_fd_sc_hd__and3_2 _09049_ (.A(_03241_),
    .B(_03250_),
    .C(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__a21oi_2 _09050_ (.A1(_03250_),
    .A2(_03251_),
    .B1(_03241_),
    .Y(_03253_));
 sky130_fd_sc_hd__a211oi_4 _09051_ (.A1(_03132_),
    .A2(_03134_),
    .B1(_03252_),
    .C1(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__o211a_1 _09052_ (.A1(_03252_),
    .A2(_03253_),
    .B1(_03132_),
    .C1(_03134_),
    .X(_03255_));
 sky130_fd_sc_hd__a211o_1 _09053_ (.A1(_03137_),
    .A2(_03139_),
    .B1(_03254_),
    .C1(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__o211ai_2 _09054_ (.A1(_03254_),
    .A2(_03255_),
    .B1(_03137_),
    .C1(_03139_),
    .Y(_03257_));
 sky130_fd_sc_hd__and3_2 _09055_ (.A(_03240_),
    .B(_03256_),
    .C(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__inv_2 _09056_ (.A(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__a21oi_2 _09057_ (.A1(_03256_),
    .A2(_03257_),
    .B1(_03240_),
    .Y(_03260_));
 sky130_fd_sc_hd__a211oi_4 _09058_ (.A1(_03141_),
    .A2(_03144_),
    .B1(_03258_),
    .C1(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__o211a_1 _09059_ (.A1(_03258_),
    .A2(_03260_),
    .B1(_03141_),
    .C1(_03144_),
    .X(_03262_));
 sky130_fd_sc_hd__nor3b_2 _09060_ (.A(_03261_),
    .B(_03262_),
    .C_N(_03224_),
    .Y(_03263_));
 sky130_fd_sc_hd__o21ba_1 _09061_ (.A1(_03261_),
    .A2(_03262_),
    .B1_N(_03224_),
    .X(_03264_));
 sky130_fd_sc_hd__a211o_1 _09062_ (.A1(_03146_),
    .A2(_03148_),
    .B1(_03263_),
    .C1(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__o211ai_2 _09063_ (.A1(_03263_),
    .A2(_03264_),
    .B1(_03146_),
    .C1(_03148_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand3b_2 _09064_ (.A_N(_03150_),
    .B(_03265_),
    .C(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__inv_2 _09065_ (.A(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21bo_1 _09066_ (.A1(_03265_),
    .A2(_03266_),
    .B1_N(_03150_),
    .X(_03269_));
 sky130_fd_sc_hd__o211a_1 _09067_ (.A1(_03120_),
    .A2(_03123_),
    .B1(_03267_),
    .C1(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__a211oi_1 _09068_ (.A1(_03267_),
    .A2(_03269_),
    .B1(_03120_),
    .C1(_03123_),
    .Y(_03271_));
 sky130_fd_sc_hd__nor2_2 _09069_ (.A(_03270_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__nand2_1 _09070_ (.A(_03200_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__xor2_2 _09071_ (.A(_03200_),
    .B(_03272_),
    .X(_03274_));
 sky130_fd_sc_hd__a21oi_1 _09072_ (.A1(_03159_),
    .A2(_03160_),
    .B1(_03158_),
    .Y(_03275_));
 sky130_fd_sc_hd__xnor2_1 _09073_ (.A(_03274_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__mux2_1 _09074_ (.A0(net3657),
    .A1(_03276_),
    .S(net484),
    .X(_03277_));
 sky130_fd_sc_hd__and3_1 _09075_ (.A(_01895_),
    .B(_01910_),
    .C(_03163_),
    .X(_03278_));
 sky130_fd_sc_hd__a21o_1 _09076_ (.A1(_01895_),
    .A2(_03163_),
    .B1(_01910_),
    .X(_03279_));
 sky130_fd_sc_hd__nand2_1 _09077_ (.A(net467),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__o2bb2a_4 _09078_ (.A1_N(net469),
    .A2_N(_03277_),
    .B1(_03278_),
    .B2(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__inv_2 _09079_ (.A(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__a21o_4 _09080_ (.A1(net391),
    .A2(_03282_),
    .B1(_03199_),
    .X(_03283_));
 sky130_fd_sc_hd__a21o_1 _09081_ (.A1(net3464),
    .A2(_01836_),
    .B1(_02946_),
    .X(_03284_));
 sky130_fd_sc_hd__and2_1 _09082_ (.A(net3241),
    .B(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__or2_1 _09083_ (.A(net3241),
    .B(_03284_),
    .X(_03286_));
 sky130_fd_sc_hd__and2b_1 _09084_ (.A_N(_03285_),
    .B(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__a21o_1 _09085_ (.A1(_03170_),
    .A2(_03172_),
    .B1(_03169_),
    .X(_03288_));
 sky130_fd_sc_hd__xnor2_1 _09086_ (.A(_03287_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__and3_1 _09087_ (.A(net3510),
    .B(net3555),
    .C(_03061_),
    .X(_03290_));
 sky130_fd_sc_hd__a21oi_1 _09088_ (.A1(net233),
    .A2(_03061_),
    .B1(net3510),
    .Y(_03291_));
 sky130_fd_sc_hd__or3_1 _09089_ (.A(_01958_),
    .B(_03290_),
    .C(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__a21oi_1 _09090_ (.A1(\dpath.btarg_DX.q[15] ),
    .A2(net403),
    .B1(net449),
    .Y(_03293_));
 sky130_fd_sc_hd__o211a_1 _09091_ (.A1(net365),
    .A2(_03289_),
    .B1(_03292_),
    .C1(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__a21bo_1 _09092_ (.A1(_02027_),
    .A2(_03283_),
    .B1_N(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__o211a_1 _09093_ (.A1(net3510),
    .A2(net441),
    .B1(_03295_),
    .C1(net845),
    .X(_00651_));
 sky130_fd_sc_hd__xnor2_1 _09094_ (.A(net3558),
    .B(_03290_),
    .Y(_03296_));
 sky130_fd_sc_hd__mux4_1 _09095_ (.A0(\dpath.RF.R[0][16] ),
    .A1(\dpath.RF.R[1][16] ),
    .A2(\dpath.RF.R[2][16] ),
    .A3(\dpath.RF.R[3][16] ),
    .S0(net567),
    .S1(net548),
    .X(_03297_));
 sky130_fd_sc_hd__mux4_1 _09096_ (.A0(\dpath.RF.R[4][16] ),
    .A1(\dpath.RF.R[5][16] ),
    .A2(\dpath.RF.R[6][16] ),
    .A3(\dpath.RF.R[7][16] ),
    .S0(net567),
    .S1(net548),
    .X(_03298_));
 sky130_fd_sc_hd__o21a_1 _09097_ (.A1(net514),
    .A2(_03298_),
    .B1(net507),
    .X(_03299_));
 sky130_fd_sc_hd__o21ai_1 _09098_ (.A1(net535),
    .A2(_03297_),
    .B1(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__mux4_1 _09099_ (.A0(\dpath.RF.R[12][16] ),
    .A1(\dpath.RF.R[13][16] ),
    .A2(\dpath.RF.R[14][16] ),
    .A3(\dpath.RF.R[15][16] ),
    .S0(net566),
    .S1(net547),
    .X(_03301_));
 sky130_fd_sc_hd__mux4_1 _09100_ (.A0(\dpath.RF.R[8][16] ),
    .A1(\dpath.RF.R[9][16] ),
    .A2(\dpath.RF.R[10][16] ),
    .A3(\dpath.RF.R[11][16] ),
    .S0(net566),
    .S1(net547),
    .X(_03302_));
 sky130_fd_sc_hd__or2_1 _09101_ (.A(net535),
    .B(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__o211a_1 _09102_ (.A1(net514),
    .A2(_03301_),
    .B1(_03303_),
    .C1(net525),
    .X(_03304_));
 sky130_fd_sc_hd__nor2_1 _09103_ (.A(net519),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__mux4_1 _09104_ (.A0(\dpath.RF.R[16][16] ),
    .A1(\dpath.RF.R[17][16] ),
    .A2(\dpath.RF.R[18][16] ),
    .A3(\dpath.RF.R[19][16] ),
    .S0(net566),
    .S1(net547),
    .X(_03306_));
 sky130_fd_sc_hd__nor2_1 _09105_ (.A(net535),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__mux4_1 _09106_ (.A0(\dpath.RF.R[20][16] ),
    .A1(\dpath.RF.R[21][16] ),
    .A2(\dpath.RF.R[22][16] ),
    .A3(\dpath.RF.R[23][16] ),
    .S0(net566),
    .S1(net547),
    .X(_03308_));
 sky130_fd_sc_hd__nor2_1 _09107_ (.A(net514),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__mux4_1 _09108_ (.A0(\dpath.RF.R[28][16] ),
    .A1(\dpath.RF.R[29][16] ),
    .A2(\dpath.RF.R[30][16] ),
    .A3(\dpath.RF.R[31][16] ),
    .S0(net566),
    .S1(net547),
    .X(_03310_));
 sky130_fd_sc_hd__nor2_1 _09109_ (.A(net514),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__mux4_1 _09110_ (.A0(\dpath.RF.R[24][16] ),
    .A1(\dpath.RF.R[25][16] ),
    .A2(\dpath.RF.R[26][16] ),
    .A3(\dpath.RF.R[27][16] ),
    .S0(net566),
    .S1(net547),
    .X(_03312_));
 sky130_fd_sc_hd__o21ai_1 _09111_ (.A1(net535),
    .A2(_03312_),
    .B1(net525),
    .Y(_03313_));
 sky130_fd_sc_hd__o32a_1 _09112_ (.A1(net525),
    .A2(_03307_),
    .A3(_03309_),
    .B1(_03311_),
    .B2(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__a221o_1 _09113_ (.A1(_03300_),
    .A2(_03305_),
    .B1(_03314_),
    .B2(net519),
    .C1(net483),
    .X(_03315_));
 sky130_fd_sc_hd__nor2_1 _09114_ (.A(net371),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__mux2_1 _09115_ (.A0(net3642),
    .A1(net8),
    .S(net480),
    .X(_03317_));
 sky130_fd_sc_hd__a221o_1 _09116_ (.A1(net686),
    .A2(net369),
    .B1(net367),
    .B2(_03317_),
    .C1(_03316_),
    .X(_03318_));
 sky130_fd_sc_hd__nand3_1 _09117_ (.A(_03045_),
    .B(_03159_),
    .C(_03274_),
    .Y(_03319_));
 sky130_fd_sc_hd__a21oi_1 _09118_ (.A1(_02935_),
    .A2(_03043_),
    .B1(_03044_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand3_1 _09119_ (.A(_03159_),
    .B(_03274_),
    .C(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__o21ai_1 _09120_ (.A1(_03200_),
    .A2(_03272_),
    .B1(_03158_),
    .Y(_03322_));
 sky130_fd_sc_hd__o2111a_2 _09121_ (.A1(_02939_),
    .A2(_03319_),
    .B1(_03321_),
    .C1(_03322_),
    .D1(_03273_),
    .X(_03323_));
 sky130_fd_sc_hd__a31oi_2 _09122_ (.A1(net788),
    .A2(net597),
    .A3(_03238_),
    .B1(_03237_),
    .Y(_03324_));
 sky130_fd_sc_hd__a22o_1 _09123_ (.A1(net649),
    .A2(net734),
    .B1(net732),
    .B2(net652),
    .X(_03325_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(net732),
    .B(_03202_),
    .Y(_03326_));
 sky130_fd_sc_hd__and4_1 _09125_ (.A(net645),
    .B(net736),
    .C(_03325_),
    .D(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__a22oi_2 _09126_ (.A1(net645),
    .A2(net736),
    .B1(_03325_),
    .B2(_03326_),
    .Y(_03328_));
 sky130_fd_sc_hd__nor3_1 _09127_ (.A(_03203_),
    .B(_03327_),
    .C(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__o21a_1 _09128_ (.A1(_03327_),
    .A2(_03328_),
    .B1(_03203_),
    .X(_03330_));
 sky130_fd_sc_hd__or2_1 _09129_ (.A(_03329_),
    .B(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__a22o_1 _09130_ (.A1(net621),
    .A2(net755),
    .B1(net752),
    .B2(net625),
    .X(_03332_));
 sky130_fd_sc_hd__and3_1 _09131_ (.A(net625),
    .B(net621),
    .C(net752),
    .X(_03333_));
 sky130_fd_sc_hd__a21bo_1 _09132_ (.A1(net755),
    .A2(_03333_),
    .B1_N(_03332_),
    .X(_03334_));
 sky130_fd_sc_hd__xor2_1 _09133_ (.A(_01864_),
    .B(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__a22o_1 _09134_ (.A1(net632),
    .A2(net745),
    .B1(net740),
    .B2(net637),
    .X(_03336_));
 sky130_fd_sc_hd__and4_1 _09135_ (.A(net637),
    .B(net633),
    .C(net744),
    .D(net740),
    .X(_03337_));
 sky130_fd_sc_hd__nand4_1 _09136_ (.A(net637),
    .B(net633),
    .C(net745),
    .D(net741),
    .Y(_03338_));
 sky130_fd_sc_hd__and4_1 _09137_ (.A(net628),
    .B(net749),
    .C(_03336_),
    .D(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__nand4_1 _09138_ (.A(net628),
    .B(net749),
    .C(_03336_),
    .D(_03338_),
    .Y(_03340_));
 sky130_fd_sc_hd__a22o_1 _09139_ (.A1(net628),
    .A2(net748),
    .B1(_03336_),
    .B2(_03338_),
    .X(_03341_));
 sky130_fd_sc_hd__o211a_1 _09140_ (.A1(_03211_),
    .A2(_03213_),
    .B1(_03340_),
    .C1(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__a211o_1 _09141_ (.A1(_03340_),
    .A2(_03341_),
    .B1(_03211_),
    .C1(_03213_),
    .X(_03343_));
 sky130_fd_sc_hd__and2b_1 _09142_ (.A_N(_03342_),
    .B(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__xnor2_1 _09143_ (.A(_03335_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__nor2_1 _09144_ (.A(_03331_),
    .B(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__and2_1 _09145_ (.A(_03331_),
    .B(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__or3_2 _09146_ (.A(_03220_),
    .B(_03346_),
    .C(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__o21ai_1 _09147_ (.A1(_03346_),
    .A2(_03347_),
    .B1(_03220_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(_03348_),
    .B(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__o21ba_1 _09149_ (.A1(_03226_),
    .A2(_03234_),
    .B1_N(_03233_),
    .X(_03351_));
 sky130_fd_sc_hd__nand2_1 _09150_ (.A(net785),
    .B(net597),
    .Y(_03352_));
 sky130_fd_sc_hd__and2_1 _09151_ (.A(net781),
    .B(net600),
    .X(_03353_));
 sky130_fd_sc_hd__a22o_1 _09152_ (.A1(net775),
    .A2(net606),
    .B1(\dpath.alu.adder.in0[13] ),
    .B2(net779),
    .X(_03354_));
 sky130_fd_sc_hd__nand4_1 _09153_ (.A(net778),
    .B(net775),
    .C(net606),
    .D(\dpath.alu.adder.in0[13] ),
    .Y(_03355_));
 sky130_fd_sc_hd__nand3_1 _09154_ (.A(_03353_),
    .B(_03354_),
    .C(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21o_1 _09155_ (.A1(_03354_),
    .A2(_03355_),
    .B1(_03353_),
    .X(_03357_));
 sky130_fd_sc_hd__a21bo_1 _09156_ (.A1(_03227_),
    .A2(_03228_),
    .B1_N(_03229_),
    .X(_03358_));
 sky130_fd_sc_hd__and3_1 _09157_ (.A(_03356_),
    .B(_03357_),
    .C(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__a21oi_1 _09158_ (.A1(_03356_),
    .A2(_03357_),
    .B1(_03358_),
    .Y(_03360_));
 sky130_fd_sc_hd__nor2_1 _09159_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xnor2_2 _09160_ (.A(_03352_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2b_1 _09161_ (.A_N(_03351_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__xnor2_2 _09162_ (.A(_03351_),
    .B(_03362_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand2_1 _09163_ (.A(net788),
    .B(net594),
    .Y(_03365_));
 sky130_fd_sc_hd__nand3_2 _09164_ (.A(net788),
    .B(net594),
    .C(_03364_),
    .Y(_03366_));
 sky130_fd_sc_hd__xnor2_1 _09165_ (.A(_03364_),
    .B(_03365_),
    .Y(_03367_));
 sky130_fd_sc_hd__a21o_1 _09166_ (.A1(_03209_),
    .A2(_03217_),
    .B1(_03216_),
    .X(_03368_));
 sky130_fd_sc_hd__nand2_1 _09167_ (.A(_03245_),
    .B(_03246_),
    .Y(_03369_));
 sky130_fd_sc_hd__a32o_1 _09168_ (.A1(net621),
    .A2(net758),
    .A3(_03206_),
    .B1(_03207_),
    .B2(net755),
    .X(_03370_));
 sky130_fd_sc_hd__a22o_1 _09169_ (.A1(net761),
    .A2(net613),
    .B1(net611),
    .B2(net766),
    .X(_03371_));
 sky130_fd_sc_hd__nand4_4 _09170_ (.A(net766),
    .B(net761),
    .C(net613),
    .D(net611),
    .Y(_03372_));
 sky130_fd_sc_hd__nand4_4 _09171_ (.A(net769),
    .B(net608),
    .C(_03371_),
    .D(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__a22o_1 _09172_ (.A1(net769),
    .A2(net608),
    .B1(_03371_),
    .B2(_03372_),
    .X(_03374_));
 sky130_fd_sc_hd__nand3_4 _09173_ (.A(_03370_),
    .B(_03373_),
    .C(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__a21o_1 _09174_ (.A1(_03373_),
    .A2(_03374_),
    .B1(_03370_),
    .X(_03376_));
 sky130_fd_sc_hd__nand3_4 _09175_ (.A(_03369_),
    .B(_03375_),
    .C(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__a21o_1 _09176_ (.A1(_03375_),
    .A2(_03376_),
    .B1(_03369_),
    .X(_03378_));
 sky130_fd_sc_hd__and3_1 _09177_ (.A(_03368_),
    .B(_03377_),
    .C(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__nand3_1 _09178_ (.A(_03368_),
    .B(_03377_),
    .C(_03378_),
    .Y(_03380_));
 sky130_fd_sc_hd__a21oi_2 _09179_ (.A1(_03377_),
    .A2(_03378_),
    .B1(_03368_),
    .Y(_03381_));
 sky130_fd_sc_hd__a211o_2 _09180_ (.A1(_03248_),
    .A2(_03250_),
    .B1(_03379_),
    .C1(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__o211ai_4 _09181_ (.A1(_03379_),
    .A2(_03381_),
    .B1(_03248_),
    .C1(_03250_),
    .Y(_03383_));
 sky130_fd_sc_hd__o211ai_4 _09182_ (.A1(_03252_),
    .A2(_03254_),
    .B1(_03382_),
    .C1(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__a211o_1 _09183_ (.A1(_03382_),
    .A2(_03383_),
    .B1(_03252_),
    .C1(_03254_),
    .X(_03385_));
 sky130_fd_sc_hd__nand3_2 _09184_ (.A(_03367_),
    .B(_03384_),
    .C(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__a21o_1 _09185_ (.A1(_03384_),
    .A2(_03385_),
    .B1(_03367_),
    .X(_03387_));
 sky130_fd_sc_hd__and3_1 _09186_ (.A(_03223_),
    .B(_03386_),
    .C(_03387_),
    .X(_03388_));
 sky130_fd_sc_hd__a21oi_1 _09187_ (.A1(_03386_),
    .A2(_03387_),
    .B1(_03223_),
    .Y(_03389_));
 sky130_fd_sc_hd__a211oi_2 _09188_ (.A1(_03256_),
    .A2(_03259_),
    .B1(_03388_),
    .C1(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__o211a_1 _09189_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03256_),
    .C1(_03259_),
    .X(_03391_));
 sky130_fd_sc_hd__or3_2 _09190_ (.A(_03350_),
    .B(_03390_),
    .C(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__o21ai_1 _09191_ (.A1(_03390_),
    .A2(_03391_),
    .B1(_03350_),
    .Y(_03393_));
 sky130_fd_sc_hd__o211ai_2 _09192_ (.A1(_03261_),
    .A2(_03263_),
    .B1(_03392_),
    .C1(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__a211o_1 _09193_ (.A1(_03392_),
    .A2(_03393_),
    .B1(_03261_),
    .C1(_03263_),
    .X(_03395_));
 sky130_fd_sc_hd__and2_1 _09194_ (.A(_03394_),
    .B(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__nand2b_1 _09195_ (.A_N(_03265_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__xnor2_1 _09196_ (.A(_03265_),
    .B(_03396_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2b_1 _09197_ (.A_N(_03324_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__xnor2_1 _09198_ (.A(_03324_),
    .B(_03398_),
    .Y(_03400_));
 sky130_fd_sc_hd__or2_1 _09199_ (.A(_03268_),
    .B(_03270_),
    .X(_03401_));
 sky130_fd_sc_hd__nand2_1 _09200_ (.A(_03400_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__or2_1 _09201_ (.A(_03400_),
    .B(_03401_),
    .X(_03403_));
 sky130_fd_sc_hd__nand2_2 _09202_ (.A(_03402_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(_03323_),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__or2_1 _09204_ (.A(_03323_),
    .B(_03404_),
    .X(_03406_));
 sky130_fd_sc_hd__nand3_1 _09205_ (.A(_01891_),
    .B(_01908_),
    .C(_03279_),
    .Y(_03407_));
 sky130_fd_sc_hd__a21o_1 _09206_ (.A1(_01908_),
    .A2(_03279_),
    .B1(_01891_),
    .X(_03408_));
 sky130_fd_sc_hd__a32o_1 _09207_ (.A1(net467),
    .A2(_03407_),
    .A3(_03408_),
    .B1(net485),
    .B2(net3453),
    .X(_03409_));
 sky130_fd_sc_hd__a31oi_4 _09208_ (.A1(_02239_),
    .A2(_03405_),
    .A3(_03406_),
    .B1(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__inv_2 _09209_ (.A(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__a21oi_4 _09210_ (.A1(net391),
    .A2(_03411_),
    .B1(_03318_),
    .Y(_03412_));
 sky130_fd_sc_hd__a21o_1 _09211_ (.A1(_03286_),
    .A2(_03288_),
    .B1(_03285_),
    .X(_03413_));
 sky130_fd_sc_hd__a21oi_1 _09212_ (.A1(net3226),
    .A2(_01836_),
    .B1(_02946_),
    .Y(_03414_));
 sky130_fd_sc_hd__and2b_1 _09213_ (.A_N(_03414_),
    .B(net3265),
    .X(_03415_));
 sky130_fd_sc_hd__and2b_1 _09214_ (.A_N(net3265),
    .B(_03414_),
    .X(_03416_));
 sky130_fd_sc_hd__nor2_1 _09215_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _09216_ (.A(_03413_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__or2_1 _09217_ (.A(_03413_),
    .B(_03417_),
    .X(_03419_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(_03418_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21oi_1 _09219_ (.A1(\dpath.btarg_DX.q[16] ),
    .A2(net403),
    .B1(net361),
    .Y(_03421_));
 sky130_fd_sc_hd__o221a_1 _09220_ (.A1(net373),
    .A2(_03412_),
    .B1(_03420_),
    .B2(net365),
    .C1(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__a21oi_1 _09221_ (.A1(net361),
    .A2(_03296_),
    .B1(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__or2_1 _09222_ (.A(net3558),
    .B(net441),
    .X(_03424_));
 sky130_fd_sc_hd__o211a_1 _09223_ (.A1(net449),
    .A2(_03423_),
    .B1(_03424_),
    .C1(net844),
    .X(_00652_));
 sky130_fd_sc_hd__mux4_1 _09224_ (.A0(\dpath.RF.R[0][17] ),
    .A1(\dpath.RF.R[1][17] ),
    .A2(\dpath.RF.R[2][17] ),
    .A3(\dpath.RF.R[3][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03425_));
 sky130_fd_sc_hd__mux4_1 _09225_ (.A0(\dpath.RF.R[4][17] ),
    .A1(\dpath.RF.R[5][17] ),
    .A2(\dpath.RF.R[6][17] ),
    .A3(\dpath.RF.R[7][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03426_));
 sky130_fd_sc_hd__o21a_1 _09226_ (.A1(net514),
    .A2(_03426_),
    .B1(net507),
    .X(_03427_));
 sky130_fd_sc_hd__o21ai_1 _09227_ (.A1(net535),
    .A2(_03425_),
    .B1(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__mux4_1 _09228_ (.A0(\dpath.RF.R[12][17] ),
    .A1(\dpath.RF.R[13][17] ),
    .A2(\dpath.RF.R[14][17] ),
    .A3(\dpath.RF.R[15][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03429_));
 sky130_fd_sc_hd__mux4_1 _09229_ (.A0(\dpath.RF.R[8][17] ),
    .A1(\dpath.RF.R[9][17] ),
    .A2(\dpath.RF.R[10][17] ),
    .A3(\dpath.RF.R[11][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03430_));
 sky130_fd_sc_hd__or2_1 _09230_ (.A(net535),
    .B(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__o211a_1 _09231_ (.A1(net514),
    .A2(_03429_),
    .B1(_03431_),
    .C1(net525),
    .X(_03432_));
 sky130_fd_sc_hd__nor2_1 _09232_ (.A(net519),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__mux4_1 _09233_ (.A0(\dpath.RF.R[16][17] ),
    .A1(\dpath.RF.R[17][17] ),
    .A2(\dpath.RF.R[18][17] ),
    .A3(\dpath.RF.R[19][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03434_));
 sky130_fd_sc_hd__nor2_1 _09234_ (.A(net535),
    .B(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__mux4_1 _09235_ (.A0(\dpath.RF.R[20][17] ),
    .A1(\dpath.RF.R[21][17] ),
    .A2(\dpath.RF.R[22][17] ),
    .A3(\dpath.RF.R[23][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03436_));
 sky130_fd_sc_hd__nor2_1 _09236_ (.A(net514),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__mux4_1 _09237_ (.A0(\dpath.RF.R[28][17] ),
    .A1(\dpath.RF.R[29][17] ),
    .A2(\dpath.RF.R[30][17] ),
    .A3(\dpath.RF.R[31][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03438_));
 sky130_fd_sc_hd__nor2_1 _09238_ (.A(net514),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__mux4_1 _09239_ (.A0(\dpath.RF.R[24][17] ),
    .A1(\dpath.RF.R[25][17] ),
    .A2(\dpath.RF.R[26][17] ),
    .A3(\dpath.RF.R[27][17] ),
    .S0(net566),
    .S1(net547),
    .X(_03440_));
 sky130_fd_sc_hd__o21ai_1 _09240_ (.A1(net535),
    .A2(_03440_),
    .B1(net525),
    .Y(_03441_));
 sky130_fd_sc_hd__o32a_1 _09241_ (.A1(net525),
    .A2(_03435_),
    .A3(_03437_),
    .B1(_03439_),
    .B2(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__a221o_1 _09242_ (.A1(_03428_),
    .A2(_03433_),
    .B1(_03442_),
    .B2(net519),
    .C1(net483),
    .X(_03443_));
 sky130_fd_sc_hd__nor2_1 _09243_ (.A(net371),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__mux2_1 _09244_ (.A0(net3633),
    .A1(net9),
    .S(net479),
    .X(_03445_));
 sky130_fd_sc_hd__a221o_1 _09245_ (.A1(net685),
    .A2(net369),
    .B1(net367),
    .B2(_03445_),
    .C1(_03444_),
    .X(_03446_));
 sky130_fd_sc_hd__nand2_1 _09246_ (.A(net758),
    .B(net615),
    .Y(_03447_));
 sky130_fd_sc_hd__a22o_1 _09247_ (.A1(net619),
    .A2(net755),
    .B1(net752),
    .B2(net623),
    .X(_03448_));
 sky130_fd_sc_hd__and3_1 _09248_ (.A(net623),
    .B(net619),
    .C(net752),
    .X(_03449_));
 sky130_fd_sc_hd__a21bo_1 _09249_ (.A1(net755),
    .A2(_03449_),
    .B1_N(_03448_),
    .X(_03450_));
 sky130_fd_sc_hd__xor2_1 _09250_ (.A(_03447_),
    .B(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__a22o_1 _09251_ (.A1(net629),
    .A2(net744),
    .B1(net741),
    .B2(net633),
    .X(_03452_));
 sky130_fd_sc_hd__and4_1 _09252_ (.A(net633),
    .B(net629),
    .C(net744),
    .D(net741),
    .X(_03453_));
 sky130_fd_sc_hd__nand4_1 _09253_ (.A(net633),
    .B(net629),
    .C(net745),
    .D(net741),
    .Y(_03454_));
 sky130_fd_sc_hd__and4_1 _09254_ (.A(net625),
    .B(net748),
    .C(_03452_),
    .D(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__nand4_1 _09255_ (.A(net625),
    .B(net748),
    .C(_03452_),
    .D(_03454_),
    .Y(_03456_));
 sky130_fd_sc_hd__a22o_1 _09256_ (.A1(net625),
    .A2(net749),
    .B1(_03452_),
    .B2(_03454_),
    .X(_03457_));
 sky130_fd_sc_hd__o211a_1 _09257_ (.A1(_03337_),
    .A2(_03339_),
    .B1(_03456_),
    .C1(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__a211o_1 _09258_ (.A1(_03456_),
    .A2(_03457_),
    .B1(_03337_),
    .C1(_03339_),
    .X(_03459_));
 sky130_fd_sc_hd__and2b_1 _09259_ (.A_N(_03458_),
    .B(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__xnor2_1 _09260_ (.A(_03451_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a22o_1 _09261_ (.A1(net645),
    .A2(net734),
    .B1(net732),
    .B2(net649),
    .X(_03462_));
 sky130_fd_sc_hd__and4_1 _09262_ (.A(net649),
    .B(net645),
    .C(net734),
    .D(net732),
    .X(_03463_));
 sky130_fd_sc_hd__inv_2 _09263_ (.A(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__and4_1 _09264_ (.A(net639),
    .B(net736),
    .C(_03462_),
    .D(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__a22oi_1 _09265_ (.A1(net639),
    .A2(net736),
    .B1(_03462_),
    .B2(_03464_),
    .Y(_03466_));
 sky130_fd_sc_hd__nor2_1 _09266_ (.A(_03465_),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__a21oi_1 _09267_ (.A1(net732),
    .A2(_03202_),
    .B1(_03327_),
    .Y(_03468_));
 sky130_fd_sc_hd__and2b_1 _09268_ (.A_N(_03468_),
    .B(_03467_),
    .X(_03469_));
 sky130_fd_sc_hd__xnor2_1 _09269_ (.A(_03467_),
    .B(_03468_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _09270_ (.A(_03329_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__xnor2_1 _09271_ (.A(_03329_),
    .B(_03470_),
    .Y(_03472_));
 sky130_fd_sc_hd__nor2_1 _09272_ (.A(_03461_),
    .B(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__or2_1 _09273_ (.A(_03461_),
    .B(_03472_),
    .X(_03474_));
 sky130_fd_sc_hd__and2_1 _09274_ (.A(_03461_),
    .B(_03472_),
    .X(_03475_));
 sky130_fd_sc_hd__or3b_2 _09275_ (.A(_03473_),
    .B(_03475_),
    .C_N(_03346_),
    .X(_03476_));
 sky130_fd_sc_hd__o21bai_1 _09276_ (.A1(_03473_),
    .A2(_03475_),
    .B1_N(_03346_),
    .Y(_03477_));
 sky130_fd_sc_hd__and4_1 _09277_ (.A(net653),
    .B(net731),
    .C(_03476_),
    .D(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__a22oi_1 _09278_ (.A1(net652),
    .A2(net731),
    .B1(_03476_),
    .B2(_03477_),
    .Y(_03479_));
 sky130_fd_sc_hd__nor2_1 _09279_ (.A(_03478_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__o21ba_1 _09280_ (.A1(_03352_),
    .A2(_03360_),
    .B1_N(_03359_),
    .X(_03481_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(net785),
    .B(net594),
    .Y(_03482_));
 sky130_fd_sc_hd__and2_1 _09282_ (.A(net781),
    .B(net597),
    .X(_03483_));
 sky130_fd_sc_hd__a22o_1 _09283_ (.A1(net773),
    .A2(net603),
    .B1(net600),
    .B2(net778),
    .X(_03484_));
 sky130_fd_sc_hd__nand4_1 _09284_ (.A(net778),
    .B(net773),
    .C(net603),
    .D(net600),
    .Y(_03485_));
 sky130_fd_sc_hd__nand3_1 _09285_ (.A(_03483_),
    .B(_03484_),
    .C(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__a21o_1 _09286_ (.A1(_03484_),
    .A2(_03485_),
    .B1(_03483_),
    .X(_03487_));
 sky130_fd_sc_hd__a21bo_1 _09287_ (.A1(_03353_),
    .A2(_03354_),
    .B1_N(_03355_),
    .X(_03488_));
 sky130_fd_sc_hd__and3_1 _09288_ (.A(_03486_),
    .B(_03487_),
    .C(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__a21oi_1 _09289_ (.A1(_03486_),
    .A2(_03487_),
    .B1(_03488_),
    .Y(_03490_));
 sky130_fd_sc_hd__nor2_1 _09290_ (.A(_03489_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__xnor2_2 _09291_ (.A(_03482_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__and2b_1 _09292_ (.A_N(_03481_),
    .B(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__xnor2_2 _09293_ (.A(_03481_),
    .B(_03492_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _09294_ (.A(net789),
    .B(net591),
    .Y(_03495_));
 sky130_fd_sc_hd__xnor2_2 _09295_ (.A(_03494_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__a21o_1 _09296_ (.A1(_03335_),
    .A2(_03343_),
    .B1(_03342_),
    .X(_03497_));
 sky130_fd_sc_hd__nand2_1 _09297_ (.A(_03372_),
    .B(_03373_),
    .Y(_03498_));
 sky130_fd_sc_hd__a32o_1 _09298_ (.A1(net617),
    .A2(net758),
    .A3(_03332_),
    .B1(_03333_),
    .B2(net755),
    .X(_03499_));
 sky130_fd_sc_hd__a22o_1 _09299_ (.A1(net761),
    .A2(net611),
    .B1(net608),
    .B2(net767),
    .X(_03500_));
 sky130_fd_sc_hd__nand4_4 _09300_ (.A(net767),
    .B(net763),
    .C(net611),
    .D(net608),
    .Y(_03501_));
 sky130_fd_sc_hd__nand4_4 _09301_ (.A(net769),
    .B(net606),
    .C(_03500_),
    .D(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__a22o_1 _09302_ (.A1(net769),
    .A2(net606),
    .B1(_03500_),
    .B2(_03501_),
    .X(_03503_));
 sky130_fd_sc_hd__nand3_4 _09303_ (.A(_03499_),
    .B(_03502_),
    .C(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21o_1 _09304_ (.A1(_03502_),
    .A2(_03503_),
    .B1(_03499_),
    .X(_03505_));
 sky130_fd_sc_hd__nand3_2 _09305_ (.A(_03498_),
    .B(_03504_),
    .C(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__a21o_1 _09306_ (.A1(_03504_),
    .A2(_03505_),
    .B1(_03498_),
    .X(_03507_));
 sky130_fd_sc_hd__and3_2 _09307_ (.A(_03497_),
    .B(_03506_),
    .C(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__a21oi_2 _09308_ (.A1(_03506_),
    .A2(_03507_),
    .B1(_03497_),
    .Y(_03509_));
 sky130_fd_sc_hd__a211oi_4 _09309_ (.A1(_03375_),
    .A2(_03377_),
    .B1(_03508_),
    .C1(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__o211a_1 _09310_ (.A1(_03508_),
    .A2(_03509_),
    .B1(_03375_),
    .C1(_03377_),
    .X(_03511_));
 sky130_fd_sc_hd__a211o_2 _09311_ (.A1(_03380_),
    .A2(_03382_),
    .B1(_03510_),
    .C1(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__o211ai_2 _09312_ (.A1(_03510_),
    .A2(_03511_),
    .B1(_03380_),
    .C1(_03382_),
    .Y(_03513_));
 sky130_fd_sc_hd__and3_1 _09313_ (.A(_03496_),
    .B(_03512_),
    .C(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__nand3_2 _09314_ (.A(_03496_),
    .B(_03512_),
    .C(_03513_),
    .Y(_03515_));
 sky130_fd_sc_hd__a21oi_1 _09315_ (.A1(_03512_),
    .A2(_03513_),
    .B1(_03496_),
    .Y(_03516_));
 sky130_fd_sc_hd__nor3_1 _09316_ (.A(_03348_),
    .B(_03514_),
    .C(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__or3_1 _09317_ (.A(_03348_),
    .B(_03514_),
    .C(_03516_),
    .X(_03518_));
 sky130_fd_sc_hd__o21a_1 _09318_ (.A1(_03514_),
    .A2(_03516_),
    .B1(_03348_),
    .X(_03519_));
 sky130_fd_sc_hd__a211o_1 _09319_ (.A1(_03384_),
    .A2(_03386_),
    .B1(_03517_),
    .C1(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__o211ai_1 _09320_ (.A1(_03517_),
    .A2(_03519_),
    .B1(_03384_),
    .C1(_03386_),
    .Y(_03521_));
 sky130_fd_sc_hd__and3_2 _09321_ (.A(_03480_),
    .B(_03520_),
    .C(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__a21oi_1 _09322_ (.A1(_03520_),
    .A2(_03521_),
    .B1(_03480_),
    .Y(_03523_));
 sky130_fd_sc_hd__nor3_1 _09323_ (.A(_03392_),
    .B(_03522_),
    .C(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__or3_1 _09324_ (.A(_03392_),
    .B(_03522_),
    .C(_03523_),
    .X(_03525_));
 sky130_fd_sc_hd__o21ai_1 _09325_ (.A1(_03522_),
    .A2(_03523_),
    .B1(_03392_),
    .Y(_03526_));
 sky130_fd_sc_hd__o211a_1 _09326_ (.A1(_03388_),
    .A2(_03390_),
    .B1(_03525_),
    .C1(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__a211oi_2 _09327_ (.A1(_03525_),
    .A2(_03526_),
    .B1(_03388_),
    .C1(_03390_),
    .Y(_03528_));
 sky130_fd_sc_hd__nor3_2 _09328_ (.A(_03394_),
    .B(_03527_),
    .C(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21a_1 _09329_ (.A1(_03527_),
    .A2(_03528_),
    .B1(_03394_),
    .X(_03530_));
 sky130_fd_sc_hd__a211oi_4 _09330_ (.A1(_03363_),
    .A2(_03366_),
    .B1(_03529_),
    .C1(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__o211a_1 _09331_ (.A1(_03529_),
    .A2(_03530_),
    .B1(_03363_),
    .C1(_03366_),
    .X(_03532_));
 sky130_fd_sc_hd__a211o_1 _09332_ (.A1(_03397_),
    .A2(_03399_),
    .B1(_03531_),
    .C1(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__o211a_1 _09333_ (.A1(_03531_),
    .A2(_03532_),
    .B1(_03397_),
    .C1(_03399_),
    .X(_03534_));
 sky130_fd_sc_hd__o211ai_1 _09334_ (.A1(_03531_),
    .A2(_03532_),
    .B1(_03397_),
    .C1(_03399_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _09335_ (.A(_03533_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__o21ai_1 _09336_ (.A1(_03323_),
    .A2(_03404_),
    .B1(_03402_),
    .Y(_03537_));
 sky130_fd_sc_hd__xnor2_1 _09337_ (.A(_03536_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__or2_1 _09338_ (.A(net3672),
    .B(net484),
    .X(_03539_));
 sky130_fd_sc_hd__o211a_1 _09339_ (.A1(net485),
    .A2(_03538_),
    .B1(_03539_),
    .C1(net468),
    .X(_03540_));
 sky130_fd_sc_hd__nand2_1 _09340_ (.A(_01890_),
    .B(_03408_),
    .Y(_03541_));
 sky130_fd_sc_hd__xor2_1 _09341_ (.A(_01863_),
    .B(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__a21o_4 _09342_ (.A1(_02101_),
    .A2(_03542_),
    .B1(_03540_),
    .X(_03543_));
 sky130_fd_sc_hd__a21o_4 _09343_ (.A1(net391),
    .A2(_03543_),
    .B1(_03446_),
    .X(_03544_));
 sky130_fd_sc_hd__and2_1 _09344_ (.A(net3496),
    .B(_01836_),
    .X(_03545_));
 sky130_fd_sc_hd__o21ai_1 _09345_ (.A1(_02946_),
    .A2(_03545_),
    .B1(net3221),
    .Y(_03546_));
 sky130_fd_sc_hd__or3_1 _09346_ (.A(net3221),
    .B(_02946_),
    .C(_03545_),
    .X(_03547_));
 sky130_fd_sc_hd__nand2_1 _09347_ (.A(_03546_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__a21oi_1 _09348_ (.A1(_03413_),
    .A2(_03417_),
    .B1(_03415_),
    .Y(_03549_));
 sky130_fd_sc_hd__xnor2_1 _09349_ (.A(_03548_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__and3_1 _09350_ (.A(net3544),
    .B(net3558),
    .C(_03290_),
    .X(_03551_));
 sky130_fd_sc_hd__a21oi_1 _09351_ (.A1(net235),
    .A2(_03290_),
    .B1(net3544),
    .Y(_03552_));
 sky130_fd_sc_hd__or3_1 _09352_ (.A(_01958_),
    .B(_03551_),
    .C(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _09353_ (.A1(\dpath.btarg_DX.q[17] ),
    .A2(net403),
    .B1(net449),
    .Y(_03554_));
 sky130_fd_sc_hd__o211a_1 _09354_ (.A1(net365),
    .A2(_03550_),
    .B1(_03553_),
    .C1(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__a21bo_1 _09355_ (.A1(_02027_),
    .A2(_03544_),
    .B1_N(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__o211a_1 _09356_ (.A1(net3544),
    .A2(net441),
    .B1(_03556_),
    .C1(net844),
    .X(_00653_));
 sky130_fd_sc_hd__xnor2_1 _09357_ (.A(net3575),
    .B(_03551_),
    .Y(_03557_));
 sky130_fd_sc_hd__mux4_1 _09358_ (.A0(\dpath.RF.R[0][18] ),
    .A1(\dpath.RF.R[1][18] ),
    .A2(\dpath.RF.R[2][18] ),
    .A3(\dpath.RF.R[3][18] ),
    .S0(net568),
    .S1(net549),
    .X(_03558_));
 sky130_fd_sc_hd__mux4_1 _09359_ (.A0(\dpath.RF.R[4][18] ),
    .A1(\dpath.RF.R[5][18] ),
    .A2(\dpath.RF.R[6][18] ),
    .A3(\dpath.RF.R[7][18] ),
    .S0(net568),
    .S1(net549),
    .X(_03559_));
 sky130_fd_sc_hd__o21a_1 _09360_ (.A1(net513),
    .A2(_03559_),
    .B1(net507),
    .X(_03560_));
 sky130_fd_sc_hd__o21ai_1 _09361_ (.A1(net534),
    .A2(_03558_),
    .B1(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__mux4_1 _09362_ (.A0(\dpath.RF.R[12][18] ),
    .A1(\dpath.RF.R[13][18] ),
    .A2(\dpath.RF.R[14][18] ),
    .A3(\dpath.RF.R[15][18] ),
    .S0(net568),
    .S1(net549),
    .X(_03562_));
 sky130_fd_sc_hd__mux4_1 _09363_ (.A0(\dpath.RF.R[8][18] ),
    .A1(\dpath.RF.R[9][18] ),
    .A2(\dpath.RF.R[10][18] ),
    .A3(\dpath.RF.R[11][18] ),
    .S0(net568),
    .S1(net549),
    .X(_03563_));
 sky130_fd_sc_hd__or2_1 _09364_ (.A(net534),
    .B(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__o211a_1 _09365_ (.A1(net513),
    .A2(_03562_),
    .B1(_03564_),
    .C1(net528),
    .X(_03565_));
 sky130_fd_sc_hd__nor2_1 _09366_ (.A(net519),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__mux4_1 _09367_ (.A0(\dpath.RF.R[16][18] ),
    .A1(\dpath.RF.R[17][18] ),
    .A2(\dpath.RF.R[18][18] ),
    .A3(\dpath.RF.R[19][18] ),
    .S0(net568),
    .S1(net549),
    .X(_03567_));
 sky130_fd_sc_hd__nor2_1 _09368_ (.A(net534),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__mux4_1 _09369_ (.A0(\dpath.RF.R[20][18] ),
    .A1(\dpath.RF.R[21][18] ),
    .A2(\dpath.RF.R[22][18] ),
    .A3(\dpath.RF.R[23][18] ),
    .S0(net569),
    .S1(net550),
    .X(_03569_));
 sky130_fd_sc_hd__nor2_1 _09370_ (.A(net513),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__mux4_1 _09371_ (.A0(\dpath.RF.R[28][18] ),
    .A1(\dpath.RF.R[29][18] ),
    .A2(\dpath.RF.R[30][18] ),
    .A3(\dpath.RF.R[31][18] ),
    .S0(net569),
    .S1(net550),
    .X(_03571_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(net514),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__mux4_1 _09373_ (.A0(\dpath.RF.R[24][18] ),
    .A1(\dpath.RF.R[25][18] ),
    .A2(\dpath.RF.R[26][18] ),
    .A3(\dpath.RF.R[27][18] ),
    .S0(net567),
    .S1(net548),
    .X(_03573_));
 sky130_fd_sc_hd__o21ai_1 _09374_ (.A1(net534),
    .A2(_03573_),
    .B1(net525),
    .Y(_03574_));
 sky130_fd_sc_hd__o32a_1 _09375_ (.A1(net528),
    .A2(_03568_),
    .A3(_03570_),
    .B1(_03572_),
    .B2(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__a221o_1 _09376_ (.A1(_03561_),
    .A2(_03566_),
    .B1(_03575_),
    .B2(net519),
    .C1(net483),
    .X(_03576_));
 sky130_fd_sc_hd__nor2_1 _09377_ (.A(net371),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__mux2_1 _09378_ (.A0(net3598),
    .A1(net10),
    .S(net479),
    .X(_03578_));
 sky130_fd_sc_hd__a221o_2 _09379_ (.A1(net682),
    .A2(net369),
    .B1(net367),
    .B2(_03578_),
    .C1(_03577_),
    .X(_03579_));
 sky130_fd_sc_hd__a31o_1 _09380_ (.A1(net789),
    .A2(net591),
    .A3(_03494_),
    .B1(_03493_),
    .X(_03580_));
 sky130_fd_sc_hd__inv_2 _09381_ (.A(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__o21ba_1 _09382_ (.A1(_03482_),
    .A2(_03490_),
    .B1_N(_03489_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2_1 _09383_ (.A(net785),
    .B(net591),
    .Y(_03583_));
 sky130_fd_sc_hd__and2_1 _09384_ (.A(net781),
    .B(net594),
    .X(_03584_));
 sky130_fd_sc_hd__a22o_1 _09385_ (.A1(net773),
    .A2(net600),
    .B1(net597),
    .B2(net778),
    .X(_03585_));
 sky130_fd_sc_hd__nand4_1 _09386_ (.A(net778),
    .B(net773),
    .C(net600),
    .D(net597),
    .Y(_03586_));
 sky130_fd_sc_hd__nand3_1 _09387_ (.A(_03584_),
    .B(_03585_),
    .C(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__a21o_1 _09388_ (.A1(_03585_),
    .A2(_03586_),
    .B1(_03584_),
    .X(_03588_));
 sky130_fd_sc_hd__a21bo_1 _09389_ (.A1(_03483_),
    .A2(_03484_),
    .B1_N(_03485_),
    .X(_03589_));
 sky130_fd_sc_hd__and3_1 _09390_ (.A(_03587_),
    .B(_03588_),
    .C(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__a21oi_1 _09391_ (.A1(_03587_),
    .A2(_03588_),
    .B1(_03589_),
    .Y(_03591_));
 sky130_fd_sc_hd__nor2_1 _09392_ (.A(_03590_),
    .B(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__xnor2_1 _09393_ (.A(_03583_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__and2b_1 _09394_ (.A_N(_03582_),
    .B(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__xnor2_1 _09395_ (.A(_03582_),
    .B(_03593_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand2_1 _09396_ (.A(net789),
    .B(net588),
    .Y(_03596_));
 sky130_fd_sc_hd__and3_1 _09397_ (.A(net789),
    .B(net588),
    .C(_03595_),
    .X(_03597_));
 sky130_fd_sc_hd__xnor2_1 _09398_ (.A(_03595_),
    .B(_03596_),
    .Y(_03598_));
 sky130_fd_sc_hd__a21o_1 _09399_ (.A1(_03451_),
    .A2(_03459_),
    .B1(_03458_),
    .X(_03599_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(_03501_),
    .B(_03502_),
    .Y(_03600_));
 sky130_fd_sc_hd__a32o_1 _09401_ (.A1(net758),
    .A2(net615),
    .A3(_03448_),
    .B1(_03449_),
    .B2(net755),
    .X(_03601_));
 sky130_fd_sc_hd__a22o_1 _09402_ (.A1(net761),
    .A2(net609),
    .B1(\dpath.alu.adder.in0[12] ),
    .B2(net766),
    .X(_03602_));
 sky130_fd_sc_hd__nand4_2 _09403_ (.A(net767),
    .B(net761),
    .C(net609),
    .D(net606),
    .Y(_03603_));
 sky130_fd_sc_hd__nand4_2 _09404_ (.A(net769),
    .B(net603),
    .C(_03602_),
    .D(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__a22o_1 _09405_ (.A1(net769),
    .A2(net603),
    .B1(_03602_),
    .B2(_03603_),
    .X(_03605_));
 sky130_fd_sc_hd__nand3_4 _09406_ (.A(_03601_),
    .B(_03604_),
    .C(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__a21o_1 _09407_ (.A1(_03604_),
    .A2(_03605_),
    .B1(_03601_),
    .X(_03607_));
 sky130_fd_sc_hd__nand3_4 _09408_ (.A(_03600_),
    .B(_03606_),
    .C(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__a21o_1 _09409_ (.A1(_03606_),
    .A2(_03607_),
    .B1(_03600_),
    .X(_03609_));
 sky130_fd_sc_hd__and3_1 _09410_ (.A(_03599_),
    .B(_03608_),
    .C(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__nand3_1 _09411_ (.A(_03599_),
    .B(_03608_),
    .C(_03609_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21oi_2 _09412_ (.A1(_03608_),
    .A2(_03609_),
    .B1(_03599_),
    .Y(_03612_));
 sky130_fd_sc_hd__a211o_2 _09413_ (.A1(_03504_),
    .A2(_03506_),
    .B1(_03610_),
    .C1(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__o211ai_4 _09414_ (.A1(_03610_),
    .A2(_03612_),
    .B1(_03504_),
    .C1(_03506_),
    .Y(_03614_));
 sky130_fd_sc_hd__o211ai_4 _09415_ (.A1(_03508_),
    .A2(_03510_),
    .B1(_03613_),
    .C1(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__a211o_1 _09416_ (.A1(_03613_),
    .A2(_03614_),
    .B1(_03508_),
    .C1(_03510_),
    .X(_03616_));
 sky130_fd_sc_hd__and3_1 _09417_ (.A(_03598_),
    .B(_03615_),
    .C(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__inv_2 _09418_ (.A(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__a21oi_1 _09419_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_03598_),
    .Y(_03619_));
 sky130_fd_sc_hd__nor3_2 _09420_ (.A(_03476_),
    .B(_03617_),
    .C(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__inv_2 _09421_ (.A(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__o21a_1 _09422_ (.A1(_03617_),
    .A2(_03619_),
    .B1(_03476_),
    .X(_03622_));
 sky130_fd_sc_hd__a211o_2 _09423_ (.A1(_03512_),
    .A2(_03515_),
    .B1(_03620_),
    .C1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__o211ai_4 _09424_ (.A1(_03620_),
    .A2(_03622_),
    .B1(_03512_),
    .C1(_03515_),
    .Y(_03624_));
 sky130_fd_sc_hd__a22oi_4 _09425_ (.A1(net649),
    .A2(net731),
    .B1(net729),
    .B2(net652),
    .Y(_03625_));
 sky130_fd_sc_hd__and3_1 _09426_ (.A(net653),
    .B(net649),
    .C(net729),
    .X(_03626_));
 sky130_fd_sc_hd__and2_2 _09427_ (.A(net731),
    .B(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(net758),
    .B(net612),
    .Y(_03628_));
 sky130_fd_sc_hd__a22o_1 _09429_ (.A1(net615),
    .A2(\dpath.alu.adder.in1[9] ),
    .B1(net751),
    .B2(net619),
    .X(_03629_));
 sky130_fd_sc_hd__and3_1 _09430_ (.A(net615),
    .B(net756),
    .C(net752),
    .X(_03630_));
 sky130_fd_sc_hd__a21bo_1 _09431_ (.A1(net619),
    .A2(_03630_),
    .B1_N(_03629_),
    .X(_03631_));
 sky130_fd_sc_hd__xor2_1 _09432_ (.A(_03628_),
    .B(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__a22o_1 _09433_ (.A1(net627),
    .A2(net744),
    .B1(net740),
    .B2(net629),
    .X(_03633_));
 sky130_fd_sc_hd__and4_1 _09434_ (.A(net629),
    .B(net625),
    .C(net745),
    .D(net741),
    .X(_03634_));
 sky130_fd_sc_hd__nand4_2 _09435_ (.A(net629),
    .B(net625),
    .C(net745),
    .D(net740),
    .Y(_03635_));
 sky130_fd_sc_hd__and4_1 _09436_ (.A(net621),
    .B(net749),
    .C(_03633_),
    .D(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__nand4_1 _09437_ (.A(net620),
    .B(net749),
    .C(_03633_),
    .D(_03635_),
    .Y(_03637_));
 sky130_fd_sc_hd__a22o_1 _09438_ (.A1(net621),
    .A2(net749),
    .B1(_03633_),
    .B2(_03635_),
    .X(_03638_));
 sky130_fd_sc_hd__o211a_1 _09439_ (.A1(_03453_),
    .A2(_03455_),
    .B1(_03637_),
    .C1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a211o_1 _09440_ (.A1(_03637_),
    .A2(_03638_),
    .B1(_03453_),
    .C1(_03455_),
    .X(_03640_));
 sky130_fd_sc_hd__and2b_1 _09441_ (.A_N(_03639_),
    .B(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__xnor2_1 _09442_ (.A(_03632_),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__a22o_1 _09443_ (.A1(net639),
    .A2(net734),
    .B1(net732),
    .B2(net645),
    .X(_03643_));
 sky130_fd_sc_hd__nand4_2 _09444_ (.A(net645),
    .B(net639),
    .C(net734),
    .D(net732),
    .Y(_03644_));
 sky130_fd_sc_hd__nand4_1 _09445_ (.A(net635),
    .B(net736),
    .C(_03643_),
    .D(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__a22o_1 _09446_ (.A1(net635),
    .A2(net736),
    .B1(_03643_),
    .B2(_03644_),
    .X(_03646_));
 sky130_fd_sc_hd__and2_1 _09447_ (.A(_03645_),
    .B(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__o21a_1 _09448_ (.A1(_03463_),
    .A2(_03465_),
    .B1(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__nor3_1 _09449_ (.A(_03463_),
    .B(_03465_),
    .C(_03647_),
    .Y(_03649_));
 sky130_fd_sc_hd__nor2_1 _09450_ (.A(_03648_),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__and2_1 _09451_ (.A(_03469_),
    .B(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__xnor2_1 _09452_ (.A(_03469_),
    .B(_03650_),
    .Y(_03652_));
 sky130_fd_sc_hd__nor2_2 _09453_ (.A(_03642_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__and2_1 _09454_ (.A(_03642_),
    .B(_03652_),
    .X(_03654_));
 sky130_fd_sc_hd__a211oi_4 _09455_ (.A1(_03471_),
    .A2(_03474_),
    .B1(_03653_),
    .C1(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o211a_1 _09456_ (.A1(_03653_),
    .A2(_03654_),
    .B1(_03471_),
    .C1(_03474_),
    .X(_03656_));
 sky130_fd_sc_hd__or4_4 _09457_ (.A(_03625_),
    .B(_03627_),
    .C(_03655_),
    .D(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__o22ai_4 _09458_ (.A1(_03625_),
    .A2(_03627_),
    .B1(_03655_),
    .B2(_03656_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand3_4 _09459_ (.A(_03478_),
    .B(_03657_),
    .C(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__a21o_1 _09460_ (.A1(_03657_),
    .A2(_03658_),
    .B1(_03478_),
    .X(_03660_));
 sky130_fd_sc_hd__nand4_4 _09461_ (.A(_03623_),
    .B(_03624_),
    .C(_03659_),
    .D(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__a22o_1 _09462_ (.A1(_03623_),
    .A2(_03624_),
    .B1(_03659_),
    .B2(_03660_),
    .X(_03662_));
 sky130_fd_sc_hd__and3_1 _09463_ (.A(_03522_),
    .B(_03661_),
    .C(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__nand3_2 _09464_ (.A(_03522_),
    .B(_03661_),
    .C(_03662_),
    .Y(_03664_));
 sky130_fd_sc_hd__a21oi_1 _09465_ (.A1(_03661_),
    .A2(_03662_),
    .B1(_03522_),
    .Y(_03665_));
 sky130_fd_sc_hd__a211o_2 _09466_ (.A1(_03518_),
    .A2(_03520_),
    .B1(_03663_),
    .C1(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__o211ai_2 _09467_ (.A1(_03663_),
    .A2(_03665_),
    .B1(_03518_),
    .C1(_03520_),
    .Y(_03667_));
 sky130_fd_sc_hd__o211a_1 _09468_ (.A1(_03524_),
    .A2(_03527_),
    .B1(_03666_),
    .C1(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__a211oi_2 _09469_ (.A1(_03666_),
    .A2(_03667_),
    .B1(_03524_),
    .C1(_03527_),
    .Y(_03669_));
 sky130_fd_sc_hd__nor3_1 _09470_ (.A(_03581_),
    .B(_03668_),
    .C(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__or3_1 _09471_ (.A(_03581_),
    .B(_03668_),
    .C(_03669_),
    .X(_03671_));
 sky130_fd_sc_hd__o21ai_1 _09472_ (.A1(_03668_),
    .A2(_03669_),
    .B1(_03581_),
    .Y(_03672_));
 sky130_fd_sc_hd__o211a_1 _09473_ (.A1(_03529_),
    .A2(_03531_),
    .B1(_03671_),
    .C1(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__a211oi_1 _09474_ (.A1(_03671_),
    .A2(_03672_),
    .B1(_03529_),
    .C1(_03531_),
    .Y(_03674_));
 sky130_fd_sc_hd__or2_1 _09475_ (.A(_03673_),
    .B(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__a21o_1 _09476_ (.A1(_03402_),
    .A2(_03533_),
    .B1(_03534_),
    .X(_03676_));
 sky130_fd_sc_hd__o31a_1 _09477_ (.A1(_03323_),
    .A2(_03404_),
    .A3(_03536_),
    .B1(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_03675_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__a21o_1 _09479_ (.A1(_03675_),
    .A2(_03677_),
    .B1(_02240_),
    .X(_03679_));
 sky130_fd_sc_hd__a31o_1 _09480_ (.A1(_01862_),
    .A2(_01890_),
    .A3(_03408_),
    .B1(_01861_),
    .X(_03680_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(_01932_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__a311o_1 _09482_ (.A1(_01862_),
    .A2(_01890_),
    .A3(_03408_),
    .B1(_01932_),
    .C1(_01861_),
    .X(_03682_));
 sky130_fd_sc_hd__a32o_1 _09483_ (.A1(net467),
    .A2(_03681_),
    .A3(_03682_),
    .B1(net485),
    .B2(net3690),
    .X(_03683_));
 sky130_fd_sc_hd__o21bai_4 _09484_ (.A1(_03678_),
    .A2(_03679_),
    .B1_N(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__a21oi_4 _09485_ (.A1(net391),
    .A2(_03684_),
    .B1(_03579_),
    .Y(_03685_));
 sky130_fd_sc_hd__a21oi_2 _09486_ (.A1(net3536),
    .A2(_01836_),
    .B1(_02946_),
    .Y(_03686_));
 sky130_fd_sc_hd__xnor2_2 _09487_ (.A(_01762_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__a21boi_1 _09488_ (.A1(_03415_),
    .A2(_03547_),
    .B1_N(_03546_),
    .Y(_03688_));
 sky130_fd_sc_hd__o21ai_1 _09489_ (.A1(_03418_),
    .A2(_03548_),
    .B1(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2b_1 _09490_ (.A_N(_03687_),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__xor2_1 _09491_ (.A(_03687_),
    .B(_03689_),
    .X(_03691_));
 sky130_fd_sc_hd__a21oi_1 _09492_ (.A1(\dpath.btarg_DX.q[18] ),
    .A2(net403),
    .B1(net362),
    .Y(_03692_));
 sky130_fd_sc_hd__o221a_1 _09493_ (.A1(net373),
    .A2(_03685_),
    .B1(_03691_),
    .B2(net365),
    .C1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__a21oi_1 _09494_ (.A1(net361),
    .A2(_03557_),
    .B1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__or2_1 _09495_ (.A(net3575),
    .B(net443),
    .X(_03695_));
 sky130_fd_sc_hd__o211a_1 _09496_ (.A1(net451),
    .A2(_03694_),
    .B1(_03695_),
    .C1(net844),
    .X(_00654_));
 sky130_fd_sc_hd__a21oi_1 _09497_ (.A1(net237),
    .A2(_03551_),
    .B1(net3525),
    .Y(_03696_));
 sky130_fd_sc_hd__and3_1 _09498_ (.A(net3525),
    .B(net237),
    .C(_03551_),
    .X(_03697_));
 sky130_fd_sc_hd__o21a_1 _09499_ (.A1(_03696_),
    .A2(_03697_),
    .B1(net362),
    .X(_03698_));
 sky130_fd_sc_hd__mux4_1 _09500_ (.A0(\dpath.RF.R[0][19] ),
    .A1(\dpath.RF.R[1][19] ),
    .A2(\dpath.RF.R[2][19] ),
    .A3(\dpath.RF.R[3][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03699_));
 sky130_fd_sc_hd__mux4_1 _09501_ (.A0(\dpath.RF.R[4][19] ),
    .A1(\dpath.RF.R[5][19] ),
    .A2(\dpath.RF.R[6][19] ),
    .A3(\dpath.RF.R[7][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03700_));
 sky130_fd_sc_hd__o21a_1 _09502_ (.A1(net514),
    .A2(_03700_),
    .B1(net507),
    .X(_03701_));
 sky130_fd_sc_hd__o21ai_1 _09503_ (.A1(net535),
    .A2(_03699_),
    .B1(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__mux4_1 _09504_ (.A0(\dpath.RF.R[12][19] ),
    .A1(\dpath.RF.R[13][19] ),
    .A2(\dpath.RF.R[14][19] ),
    .A3(\dpath.RF.R[15][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03703_));
 sky130_fd_sc_hd__mux4_1 _09505_ (.A0(\dpath.RF.R[8][19] ),
    .A1(\dpath.RF.R[9][19] ),
    .A2(\dpath.RF.R[10][19] ),
    .A3(\dpath.RF.R[11][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03704_));
 sky130_fd_sc_hd__or2_1 _09506_ (.A(net535),
    .B(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__o211a_1 _09507_ (.A1(net514),
    .A2(_03703_),
    .B1(_03705_),
    .C1(net525),
    .X(_03706_));
 sky130_fd_sc_hd__nor2_1 _09508_ (.A(net519),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__mux4_1 _09509_ (.A0(\dpath.RF.R[16][19] ),
    .A1(\dpath.RF.R[17][19] ),
    .A2(\dpath.RF.R[18][19] ),
    .A3(\dpath.RF.R[19][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03708_));
 sky130_fd_sc_hd__nor2_1 _09510_ (.A(net535),
    .B(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__mux4_1 _09511_ (.A0(\dpath.RF.R[20][19] ),
    .A1(\dpath.RF.R[21][19] ),
    .A2(\dpath.RF.R[22][19] ),
    .A3(\dpath.RF.R[23][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03710_));
 sky130_fd_sc_hd__nor2_1 _09512_ (.A(net514),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__mux4_1 _09513_ (.A0(\dpath.RF.R[28][19] ),
    .A1(\dpath.RF.R[29][19] ),
    .A2(\dpath.RF.R[30][19] ),
    .A3(\dpath.RF.R[31][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03712_));
 sky130_fd_sc_hd__nor2_1 _09514_ (.A(net514),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__mux4_1 _09515_ (.A0(\dpath.RF.R[24][19] ),
    .A1(\dpath.RF.R[25][19] ),
    .A2(\dpath.RF.R[26][19] ),
    .A3(\dpath.RF.R[27][19] ),
    .S0(net567),
    .S1(net548),
    .X(_03714_));
 sky130_fd_sc_hd__o21ai_1 _09516_ (.A1(net535),
    .A2(_03714_),
    .B1(net525),
    .Y(_03715_));
 sky130_fd_sc_hd__o32a_1 _09517_ (.A1(net525),
    .A2(_03709_),
    .A3(_03711_),
    .B1(_03713_),
    .B2(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__a221o_1 _09518_ (.A1(_03702_),
    .A2(_03707_),
    .B1(_03716_),
    .B2(net519),
    .C1(net483),
    .X(_03717_));
 sky130_fd_sc_hd__nor2_1 _09519_ (.A(net371),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__mux2_2 _09520_ (.A0(net3606),
    .A1(net11),
    .S(net479),
    .X(_03719_));
 sky130_fd_sc_hd__a221o_2 _09521_ (.A1(net998),
    .A2(net369),
    .B1(net367),
    .B2(_03719_),
    .C1(_03718_),
    .X(_03720_));
 sky130_fd_sc_hd__o21ba_1 _09522_ (.A1(_03583_),
    .A2(_03591_),
    .B1_N(_03590_),
    .X(_03721_));
 sky130_fd_sc_hd__nand2_1 _09523_ (.A(net785),
    .B(net588),
    .Y(_03722_));
 sky130_fd_sc_hd__and2_1 _09524_ (.A(net781),
    .B(net591),
    .X(_03723_));
 sky130_fd_sc_hd__a22o_1 _09525_ (.A1(net773),
    .A2(net597),
    .B1(net594),
    .B2(net778),
    .X(_03724_));
 sky130_fd_sc_hd__nand4_1 _09526_ (.A(net778),
    .B(net773),
    .C(net597),
    .D(net594),
    .Y(_03725_));
 sky130_fd_sc_hd__nand3_1 _09527_ (.A(_03723_),
    .B(_03724_),
    .C(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__a21o_1 _09528_ (.A1(_03724_),
    .A2(_03725_),
    .B1(_03723_),
    .X(_03727_));
 sky130_fd_sc_hd__a21bo_1 _09529_ (.A1(_03584_),
    .A2(_03585_),
    .B1_N(_03586_),
    .X(_03728_));
 sky130_fd_sc_hd__and3_1 _09530_ (.A(_03726_),
    .B(_03727_),
    .C(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a21oi_1 _09531_ (.A1(_03726_),
    .A2(_03727_),
    .B1(_03728_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _09532_ (.A(_03729_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__xnor2_2 _09533_ (.A(_03722_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__and2b_1 _09534_ (.A_N(_03721_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__xnor2_2 _09535_ (.A(_03721_),
    .B(_03732_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _09536_ (.A(net789),
    .B(net586),
    .Y(_03735_));
 sky130_fd_sc_hd__xnor2_2 _09537_ (.A(_03734_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__a21o_1 _09538_ (.A1(_03632_),
    .A2(_03640_),
    .B1(_03639_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_1 _09539_ (.A(_03603_),
    .B(_03604_),
    .Y(_03738_));
 sky130_fd_sc_hd__a32o_1 _09540_ (.A1(net758),
    .A2(net612),
    .A3(_03629_),
    .B1(_03630_),
    .B2(net619),
    .X(_03739_));
 sky130_fd_sc_hd__a22o_1 _09541_ (.A1(net761),
    .A2(\dpath.alu.adder.in0[12] ),
    .B1(net603),
    .B2(net766),
    .X(_03740_));
 sky130_fd_sc_hd__nand4_2 _09542_ (.A(net767),
    .B(net761),
    .C(\dpath.alu.adder.in0[12] ),
    .D(net603),
    .Y(_03741_));
 sky130_fd_sc_hd__nand4_2 _09543_ (.A(net771),
    .B(net600),
    .C(_03740_),
    .D(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__a22o_1 _09544_ (.A1(net771),
    .A2(net600),
    .B1(_03740_),
    .B2(_03741_),
    .X(_03743_));
 sky130_fd_sc_hd__nand3_4 _09545_ (.A(_03739_),
    .B(_03742_),
    .C(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__a21o_1 _09546_ (.A1(_03742_),
    .A2(_03743_),
    .B1(_03739_),
    .X(_03745_));
 sky130_fd_sc_hd__nand3_2 _09547_ (.A(_03738_),
    .B(_03744_),
    .C(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21o_1 _09548_ (.A1(_03744_),
    .A2(_03745_),
    .B1(_03738_),
    .X(_03747_));
 sky130_fd_sc_hd__and3_2 _09549_ (.A(_03737_),
    .B(_03746_),
    .C(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__a21oi_2 _09550_ (.A1(_03746_),
    .A2(_03747_),
    .B1(_03737_),
    .Y(_03749_));
 sky130_fd_sc_hd__a211oi_4 _09551_ (.A1(_03606_),
    .A2(_03608_),
    .B1(_03748_),
    .C1(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__o211a_1 _09552_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_03606_),
    .C1(_03608_),
    .X(_03751_));
 sky130_fd_sc_hd__a211o_1 _09553_ (.A1(_03611_),
    .A2(_03613_),
    .B1(_03750_),
    .C1(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__o211ai_2 _09554_ (.A1(_03750_),
    .A2(_03751_),
    .B1(_03611_),
    .C1(_03613_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand3_2 _09555_ (.A(_03736_),
    .B(_03752_),
    .C(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__a21o_1 _09556_ (.A1(_03752_),
    .A2(_03753_),
    .B1(_03736_),
    .X(_03755_));
 sky130_fd_sc_hd__and3_2 _09557_ (.A(_03655_),
    .B(_03754_),
    .C(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__a21oi_2 _09558_ (.A1(_03754_),
    .A2(_03755_),
    .B1(_03655_),
    .Y(_03757_));
 sky130_fd_sc_hd__a211oi_4 _09559_ (.A1(_03615_),
    .A2(_03618_),
    .B1(_03756_),
    .C1(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__o211a_1 _09560_ (.A1(_03756_),
    .A2(_03757_),
    .B1(_03615_),
    .C1(_03618_),
    .X(_03759_));
 sky130_fd_sc_hd__nand2_1 _09561_ (.A(net645),
    .B(net731),
    .Y(_03760_));
 sky130_fd_sc_hd__a22o_1 _09562_ (.A1(net649),
    .A2(net729),
    .B1(net727),
    .B2(net653),
    .X(_03761_));
 sky130_fd_sc_hd__a21bo_1 _09563_ (.A1(net727),
    .A2(_03626_),
    .B1_N(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__xor2_1 _09564_ (.A(_03760_),
    .B(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__nand2_1 _09565_ (.A(net758),
    .B(net609),
    .Y(_03764_));
 sky130_fd_sc_hd__a22o_1 _09566_ (.A1(net755),
    .A2(net612),
    .B1(net752),
    .B2(net615),
    .X(_03765_));
 sky130_fd_sc_hd__a21bo_1 _09567_ (.A1(net612),
    .A2(_03630_),
    .B1_N(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__xor2_1 _09568_ (.A(_03764_),
    .B(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__a22o_1 _09569_ (.A1(net621),
    .A2(net745),
    .B1(net740),
    .B2(net625),
    .X(_03768_));
 sky130_fd_sc_hd__and4_1 _09570_ (.A(net625),
    .B(net621),
    .C(net745),
    .D(net741),
    .X(_03769_));
 sky130_fd_sc_hd__nand4_2 _09571_ (.A(net625),
    .B(net621),
    .C(net745),
    .D(net740),
    .Y(_03770_));
 sky130_fd_sc_hd__and4_1 _09572_ (.A(net616),
    .B(net749),
    .C(_03768_),
    .D(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__nand4_1 _09573_ (.A(net616),
    .B(net749),
    .C(_03768_),
    .D(_03770_),
    .Y(_03772_));
 sky130_fd_sc_hd__a22o_1 _09574_ (.A1(net616),
    .A2(net749),
    .B1(_03768_),
    .B2(_03770_),
    .X(_03773_));
 sky130_fd_sc_hd__o211a_1 _09575_ (.A1(_03634_),
    .A2(_03636_),
    .B1(_03772_),
    .C1(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__a211o_1 _09576_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03634_),
    .C1(_03636_),
    .X(_03775_));
 sky130_fd_sc_hd__and2b_1 _09577_ (.A_N(_03774_),
    .B(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__xnor2_1 _09578_ (.A(_03767_),
    .B(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand2_1 _09579_ (.A(_03644_),
    .B(_03645_),
    .Y(_03778_));
 sky130_fd_sc_hd__a22o_1 _09580_ (.A1(net635),
    .A2(net734),
    .B1(net732),
    .B2(net639),
    .X(_03779_));
 sky130_fd_sc_hd__and4_1 _09581_ (.A(net639),
    .B(net635),
    .C(net734),
    .D(net732),
    .X(_03780_));
 sky130_fd_sc_hd__nand4_1 _09582_ (.A(net639),
    .B(net635),
    .C(net734),
    .D(net732),
    .Y(_03781_));
 sky130_fd_sc_hd__a22oi_1 _09583_ (.A1(net631),
    .A2(net736),
    .B1(_03779_),
    .B2(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__and4_1 _09584_ (.A(net631),
    .B(net736),
    .C(_03779_),
    .D(_03781_),
    .X(_03783_));
 sky130_fd_sc_hd__nor2_1 _09585_ (.A(_03782_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__and2_1 _09586_ (.A(_03627_),
    .B(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__xnor2_1 _09587_ (.A(_03627_),
    .B(_03784_),
    .Y(_03786_));
 sky130_fd_sc_hd__and2b_1 _09588_ (.A_N(_03786_),
    .B(_03778_),
    .X(_03787_));
 sky130_fd_sc_hd__xnor2_1 _09589_ (.A(_03778_),
    .B(_03786_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(_03648_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__xnor2_1 _09591_ (.A(_03648_),
    .B(_03788_),
    .Y(_03790_));
 sky130_fd_sc_hd__or2_2 _09592_ (.A(_03777_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__nand2_1 _09593_ (.A(_03777_),
    .B(_03790_),
    .Y(_03792_));
 sky130_fd_sc_hd__o211a_1 _09594_ (.A1(_03651_),
    .A2(_03653_),
    .B1(_03791_),
    .C1(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__o211ai_1 _09595_ (.A1(_03651_),
    .A2(_03653_),
    .B1(_03791_),
    .C1(_03792_),
    .Y(_03794_));
 sky130_fd_sc_hd__a211o_1 _09596_ (.A1(_03791_),
    .A2(_03792_),
    .B1(_03651_),
    .C1(_03653_),
    .X(_03795_));
 sky130_fd_sc_hd__and3_1 _09597_ (.A(_03763_),
    .B(_03794_),
    .C(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__a21oi_1 _09598_ (.A1(_03794_),
    .A2(_03795_),
    .B1(_03763_),
    .Y(_03797_));
 sky130_fd_sc_hd__or3_4 _09599_ (.A(_03657_),
    .B(_03796_),
    .C(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__o21ai_2 _09600_ (.A1(_03796_),
    .A2(_03797_),
    .B1(_03657_),
    .Y(_03799_));
 sky130_fd_sc_hd__and4bb_1 _09601_ (.A_N(_03758_),
    .B_N(_03759_),
    .C(_03798_),
    .D(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__or4bb_2 _09602_ (.A(_03758_),
    .B(_03759_),
    .C_N(_03798_),
    .D_N(_03799_),
    .X(_03801_));
 sky130_fd_sc_hd__a2bb2oi_2 _09603_ (.A1_N(_03758_),
    .A2_N(_03759_),
    .B1(_03798_),
    .B2(_03799_),
    .Y(_03802_));
 sky130_fd_sc_hd__a211oi_4 _09604_ (.A1(_03659_),
    .A2(_03661_),
    .B1(_03800_),
    .C1(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__o211a_1 _09605_ (.A1(_03800_),
    .A2(_03802_),
    .B1(_03659_),
    .C1(_03661_),
    .X(_03804_));
 sky130_fd_sc_hd__a211oi_4 _09606_ (.A1(_03621_),
    .A2(_03623_),
    .B1(_03803_),
    .C1(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__o211a_1 _09607_ (.A1(_03803_),
    .A2(_03804_),
    .B1(_03621_),
    .C1(_03623_),
    .X(_03806_));
 sky130_fd_sc_hd__a211o_2 _09608_ (.A1(_03664_),
    .A2(_03666_),
    .B1(_03805_),
    .C1(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__o211ai_4 _09609_ (.A1(_03805_),
    .A2(_03806_),
    .B1(_03664_),
    .C1(_03666_),
    .Y(_03808_));
 sky130_fd_sc_hd__o211ai_4 _09610_ (.A1(_03594_),
    .A2(_03597_),
    .B1(_03807_),
    .C1(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__a211o_1 _09611_ (.A1(_03807_),
    .A2(_03808_),
    .B1(_03594_),
    .C1(_03597_),
    .X(_03810_));
 sky130_fd_sc_hd__a211o_1 _09612_ (.A1(_03809_),
    .A2(_03810_),
    .B1(_03668_),
    .C1(_03670_),
    .X(_03811_));
 sky130_fd_sc_hd__o211ai_2 _09613_ (.A1(_03668_),
    .A2(_03670_),
    .B1(_03809_),
    .C1(_03810_),
    .Y(_03812_));
 sky130_fd_sc_hd__nand2_1 _09614_ (.A(_03811_),
    .B(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__nor2_1 _09615_ (.A(_03673_),
    .B(_03678_),
    .Y(_03814_));
 sky130_fd_sc_hd__xor2_1 _09616_ (.A(_03813_),
    .B(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__or2_1 _09617_ (.A(net3649),
    .B(_02071_),
    .X(_03816_));
 sky130_fd_sc_hd__o211a_1 _09618_ (.A1(net486),
    .A2(_03815_),
    .B1(_03816_),
    .C1(net468),
    .X(_03817_));
 sky130_fd_sc_hd__nand3_1 _09619_ (.A(_01913_),
    .B(_01930_),
    .C(_03682_),
    .Y(_03818_));
 sky130_fd_sc_hd__a21o_1 _09620_ (.A1(_01930_),
    .A2(_03682_),
    .B1(_01913_),
    .X(_03819_));
 sky130_fd_sc_hd__a31o_4 _09621_ (.A1(_02101_),
    .A2(_03818_),
    .A3(_03819_),
    .B1(_03817_),
    .X(_03820_));
 sky130_fd_sc_hd__a21oi_4 _09622_ (.A1(net391),
    .A2(_03820_),
    .B1(_03720_),
    .Y(_03821_));
 sky130_fd_sc_hd__a21o_1 _09623_ (.A1(net3495),
    .A2(_01836_),
    .B1(_02946_),
    .X(_03822_));
 sky130_fd_sc_hd__nand2_1 _09624_ (.A(net3323),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__or2_1 _09625_ (.A(net3323),
    .B(_03822_),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_1 _09626_ (.A(_03823_),
    .B(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__o21a_1 _09627_ (.A1(_01762_),
    .A2(_03686_),
    .B1(_03690_),
    .X(_03826_));
 sky130_fd_sc_hd__xnor2_1 _09628_ (.A(_03825_),
    .B(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__a21oi_1 _09629_ (.A1(\dpath.btarg_DX.q[19] ),
    .A2(net403),
    .B1(net362),
    .Y(_03828_));
 sky130_fd_sc_hd__o221a_1 _09630_ (.A1(net373),
    .A2(_03821_),
    .B1(_03827_),
    .B2(net365),
    .C1(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__o21ai_1 _09631_ (.A1(_03698_),
    .A2(_03829_),
    .B1(net443),
    .Y(_03830_));
 sky130_fd_sc_hd__o211a_1 _09632_ (.A1(net3525),
    .A2(net443),
    .B1(_03830_),
    .C1(net844),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _09633_ (.A0(\dpath.RF.R[0][20] ),
    .A1(\dpath.RF.R[1][20] ),
    .A2(\dpath.RF.R[2][20] ),
    .A3(\dpath.RF.R[3][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03831_));
 sky130_fd_sc_hd__mux4_1 _09634_ (.A0(\dpath.RF.R[4][20] ),
    .A1(\dpath.RF.R[5][20] ),
    .A2(\dpath.RF.R[6][20] ),
    .A3(\dpath.RF.R[7][20] ),
    .S0(net570),
    .S1(net551),
    .X(_03832_));
 sky130_fd_sc_hd__o21a_1 _09635_ (.A1(net513),
    .A2(_03832_),
    .B1(net507),
    .X(_03833_));
 sky130_fd_sc_hd__o21ai_1 _09636_ (.A1(net534),
    .A2(_03831_),
    .B1(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__mux4_1 _09637_ (.A0(\dpath.RF.R[12][20] ),
    .A1(\dpath.RF.R[13][20] ),
    .A2(\dpath.RF.R[14][20] ),
    .A3(\dpath.RF.R[15][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03835_));
 sky130_fd_sc_hd__mux4_1 _09638_ (.A0(\dpath.RF.R[8][20] ),
    .A1(\dpath.RF.R[9][20] ),
    .A2(\dpath.RF.R[10][20] ),
    .A3(\dpath.RF.R[11][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03836_));
 sky130_fd_sc_hd__or2_1 _09639_ (.A(net534),
    .B(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__o211a_1 _09640_ (.A1(net513),
    .A2(_03835_),
    .B1(_03837_),
    .C1(net525),
    .X(_03838_));
 sky130_fd_sc_hd__nor2_1 _09641_ (.A(net519),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__mux4_1 _09642_ (.A0(\dpath.RF.R[16][20] ),
    .A1(\dpath.RF.R[17][20] ),
    .A2(\dpath.RF.R[18][20] ),
    .A3(\dpath.RF.R[19][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03840_));
 sky130_fd_sc_hd__nor2_1 _09643_ (.A(net534),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__mux4_1 _09644_ (.A0(\dpath.RF.R[20][20] ),
    .A1(\dpath.RF.R[21][20] ),
    .A2(\dpath.RF.R[22][20] ),
    .A3(\dpath.RF.R[23][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03842_));
 sky130_fd_sc_hd__nor2_1 _09645_ (.A(net513),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__mux4_1 _09646_ (.A0(\dpath.RF.R[28][20] ),
    .A1(\dpath.RF.R[29][20] ),
    .A2(\dpath.RF.R[30][20] ),
    .A3(\dpath.RF.R[31][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03844_));
 sky130_fd_sc_hd__nor2_1 _09647_ (.A(net513),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__mux4_1 _09648_ (.A0(\dpath.RF.R[24][20] ),
    .A1(\dpath.RF.R[25][20] ),
    .A2(\dpath.RF.R[26][20] ),
    .A3(\dpath.RF.R[27][20] ),
    .S0(net568),
    .S1(net549),
    .X(_03846_));
 sky130_fd_sc_hd__o21ai_1 _09649_ (.A1(net534),
    .A2(_03846_),
    .B1(net525),
    .Y(_03847_));
 sky130_fd_sc_hd__o32a_1 _09650_ (.A1(net525),
    .A2(_03841_),
    .A3(_03843_),
    .B1(_03845_),
    .B2(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__a221o_1 _09651_ (.A1(_03834_),
    .A2(_03839_),
    .B1(_03848_),
    .B2(net519),
    .C1(net483),
    .X(_03849_));
 sky130_fd_sc_hd__nor2_1 _09652_ (.A(net371),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(net3643),
    .A1(net13),
    .S(net479),
    .X(_03851_));
 sky130_fd_sc_hd__a221o_1 _09654_ (.A1(net679),
    .A2(net369),
    .B1(net367),
    .B2(_03851_),
    .C1(_03850_),
    .X(_03852_));
 sky130_fd_sc_hd__a31o_1 _09655_ (.A1(net789),
    .A2(net586),
    .A3(_03734_),
    .B1(_03733_),
    .X(_03853_));
 sky130_fd_sc_hd__o21ba_1 _09656_ (.A1(_03722_),
    .A2(_03730_),
    .B1_N(_03729_),
    .X(_03854_));
 sky130_fd_sc_hd__nand2_1 _09657_ (.A(net785),
    .B(net586),
    .Y(_03855_));
 sky130_fd_sc_hd__a22o_1 _09658_ (.A1(net773),
    .A2(net594),
    .B1(net591),
    .B2(net778),
    .X(_03856_));
 sky130_fd_sc_hd__nand4_2 _09659_ (.A(net778),
    .B(net773),
    .C(net594),
    .D(net591),
    .Y(_03857_));
 sky130_fd_sc_hd__a22o_1 _09660_ (.A1(net781),
    .A2(net588),
    .B1(_03856_),
    .B2(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__nand4_1 _09661_ (.A(net781),
    .B(net588),
    .C(_03856_),
    .D(_03857_),
    .Y(_03859_));
 sky130_fd_sc_hd__a21bo_1 _09662_ (.A1(_03723_),
    .A2(_03724_),
    .B1_N(_03725_),
    .X(_03860_));
 sky130_fd_sc_hd__and3_1 _09663_ (.A(_03858_),
    .B(_03859_),
    .C(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__a21oi_1 _09664_ (.A1(_03858_),
    .A2(_03859_),
    .B1(_03860_),
    .Y(_03862_));
 sky130_fd_sc_hd__nor2_1 _09665_ (.A(_03861_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__xnor2_1 _09666_ (.A(_03855_),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand2b_1 _09667_ (.A_N(_03854_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__xnor2_1 _09668_ (.A(_03854_),
    .B(_03864_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _09669_ (.A(net789),
    .B(net584),
    .Y(_03867_));
 sky130_fd_sc_hd__nand3_1 _09670_ (.A(net789),
    .B(net584),
    .C(_03866_),
    .Y(_03868_));
 sky130_fd_sc_hd__xnor2_1 _09671_ (.A(_03866_),
    .B(_03867_),
    .Y(_03869_));
 sky130_fd_sc_hd__a21o_1 _09672_ (.A1(_03767_),
    .A2(_03775_),
    .B1(_03774_),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _09673_ (.A(_03741_),
    .B(_03742_),
    .Y(_03871_));
 sky130_fd_sc_hd__a32o_1 _09674_ (.A1(net758),
    .A2(net609),
    .A3(_03765_),
    .B1(_03630_),
    .B2(net612),
    .X(_03872_));
 sky130_fd_sc_hd__a22o_1 _09675_ (.A1(net761),
    .A2(net603),
    .B1(net600),
    .B2(net766),
    .X(_03873_));
 sky130_fd_sc_hd__nand4_4 _09676_ (.A(net766),
    .B(net761),
    .C(net603),
    .D(net600),
    .Y(_03874_));
 sky130_fd_sc_hd__a22o_1 _09677_ (.A1(net769),
    .A2(net597),
    .B1(_03873_),
    .B2(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__nand4_4 _09678_ (.A(net769),
    .B(net597),
    .C(_03873_),
    .D(_03874_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand3_4 _09679_ (.A(_03872_),
    .B(_03875_),
    .C(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__a21o_1 _09680_ (.A1(_03875_),
    .A2(_03876_),
    .B1(_03872_),
    .X(_03878_));
 sky130_fd_sc_hd__nand3_4 _09681_ (.A(_03871_),
    .B(_03877_),
    .C(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__a21o_1 _09682_ (.A1(_03877_),
    .A2(_03878_),
    .B1(_03871_),
    .X(_03880_));
 sky130_fd_sc_hd__and3_1 _09683_ (.A(_03870_),
    .B(_03879_),
    .C(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__nand3_1 _09684_ (.A(_03870_),
    .B(_03879_),
    .C(_03880_),
    .Y(_03882_));
 sky130_fd_sc_hd__a21oi_2 _09685_ (.A1(_03879_),
    .A2(_03880_),
    .B1(_03870_),
    .Y(_03883_));
 sky130_fd_sc_hd__a211o_2 _09686_ (.A1(_03744_),
    .A2(_03746_),
    .B1(_03881_),
    .C1(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__o211ai_4 _09687_ (.A1(_03881_),
    .A2(_03883_),
    .B1(_03744_),
    .C1(_03746_),
    .Y(_03885_));
 sky130_fd_sc_hd__o211ai_4 _09688_ (.A1(_03748_),
    .A2(_03750_),
    .B1(_03884_),
    .C1(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__a211o_1 _09689_ (.A1(_03884_),
    .A2(_03885_),
    .B1(_03748_),
    .C1(_03750_),
    .X(_03887_));
 sky130_fd_sc_hd__nand3_2 _09690_ (.A(_03869_),
    .B(_03886_),
    .C(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__a21o_1 _09691_ (.A1(_03886_),
    .A2(_03887_),
    .B1(_03869_),
    .X(_03889_));
 sky130_fd_sc_hd__and3_1 _09692_ (.A(_03793_),
    .B(_03888_),
    .C(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__inv_2 _09693_ (.A(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__a21oi_1 _09694_ (.A1(_03888_),
    .A2(_03889_),
    .B1(_03793_),
    .Y(_03892_));
 sky130_fd_sc_hd__a211oi_2 _09695_ (.A1(_03752_),
    .A2(_03754_),
    .B1(_03890_),
    .C1(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__inv_2 _09696_ (.A(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__o211a_1 _09697_ (.A1(_03890_),
    .A2(_03892_),
    .B1(_03752_),
    .C1(_03754_),
    .X(_03895_));
 sky130_fd_sc_hd__nand2_1 _09698_ (.A(net653),
    .B(\dpath.alu.adder.in1[20] ),
    .Y(_03896_));
 sky130_fd_sc_hd__a22o_1 _09699_ (.A1(net645),
    .A2(net729),
    .B1(net727),
    .B2(net649),
    .X(_03897_));
 sky130_fd_sc_hd__inv_2 _09700_ (.A(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__and4_1 _09701_ (.A(net649),
    .B(net645),
    .C(net729),
    .D(net727),
    .X(_03899_));
 sky130_fd_sc_hd__and4b_1 _09702_ (.A_N(_03899_),
    .B(net731),
    .C(net639),
    .D(_03897_),
    .X(_03900_));
 sky130_fd_sc_hd__o2bb2a_1 _09703_ (.A1_N(net639),
    .A2_N(net731),
    .B1(_03898_),
    .B2(_03899_),
    .X(_03901_));
 sky130_fd_sc_hd__nor2_1 _09704_ (.A(_03900_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__nand2b_1 _09705_ (.A_N(_03896_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__xnor2_1 _09706_ (.A(_03896_),
    .B(_03902_),
    .Y(_03904_));
 sky130_fd_sc_hd__a22o_1 _09707_ (.A1(net612),
    .A2(net752),
    .B1(net608),
    .B2(net755),
    .X(_03905_));
 sky130_fd_sc_hd__nand4_4 _09708_ (.A(net755),
    .B(net612),
    .C(net752),
    .D(net608),
    .Y(_03906_));
 sky130_fd_sc_hd__nand4_2 _09709_ (.A(net758),
    .B(net606),
    .C(_03905_),
    .D(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__a22o_1 _09710_ (.A1(net758),
    .A2(net606),
    .B1(_03905_),
    .B2(_03906_),
    .X(_03908_));
 sky130_fd_sc_hd__and2_2 _09711_ (.A(_03907_),
    .B(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__and2_1 _09712_ (.A(net613),
    .B(net749),
    .X(_03910_));
 sky130_fd_sc_hd__a22o_1 _09713_ (.A1(net616),
    .A2(net745),
    .B1(net741),
    .B2(net621),
    .X(_03911_));
 sky130_fd_sc_hd__nand4_1 _09714_ (.A(net621),
    .B(net616),
    .C(net745),
    .D(net741),
    .Y(_03912_));
 sky130_fd_sc_hd__nand3_1 _09715_ (.A(_03910_),
    .B(_03911_),
    .C(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__a21o_1 _09716_ (.A1(_03911_),
    .A2(_03912_),
    .B1(_03910_),
    .X(_03914_));
 sky130_fd_sc_hd__o211a_1 _09717_ (.A1(_03769_),
    .A2(_03771_),
    .B1(_03913_),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__a211o_1 _09718_ (.A1(_03913_),
    .A2(_03914_),
    .B1(_03769_),
    .C1(_03771_),
    .X(_03916_));
 sky130_fd_sc_hd__and2b_1 _09719_ (.A_N(_03915_),
    .B(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__xnor2_4 _09720_ (.A(_03909_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__nor2_1 _09721_ (.A(_03780_),
    .B(_03783_),
    .Y(_03919_));
 sky130_fd_sc_hd__a32o_1 _09722_ (.A1(net645),
    .A2(net731),
    .A3(_03761_),
    .B1(_03626_),
    .B2(net727),
    .X(_03920_));
 sky130_fd_sc_hd__a22o_1 _09723_ (.A1(net631),
    .A2(net734),
    .B1(net732),
    .B2(net635),
    .X(_03921_));
 sky130_fd_sc_hd__nand4_1 _09724_ (.A(net635),
    .B(net631),
    .C(net734),
    .D(net732),
    .Y(_03922_));
 sky130_fd_sc_hd__a22oi_1 _09725_ (.A1(net627),
    .A2(net736),
    .B1(_03921_),
    .B2(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__and4_1 _09726_ (.A(net627),
    .B(net736),
    .C(_03921_),
    .D(_03922_),
    .X(_03924_));
 sky130_fd_sc_hd__or2_1 _09727_ (.A(_03923_),
    .B(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__nand2b_1 _09728_ (.A_N(_03925_),
    .B(_03920_),
    .Y(_03926_));
 sky130_fd_sc_hd__xnor2_1 _09729_ (.A(_03920_),
    .B(_03925_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2b_1 _09730_ (.A_N(_03919_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__xnor2_1 _09731_ (.A(_03919_),
    .B(_03927_),
    .Y(_03929_));
 sky130_fd_sc_hd__o21a_2 _09732_ (.A1(_03785_),
    .A2(_03787_),
    .B1(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__nor3_2 _09733_ (.A(_03785_),
    .B(_03787_),
    .C(_03929_),
    .Y(_03931_));
 sky130_fd_sc_hd__nor3_4 _09734_ (.A(_03918_),
    .B(_03930_),
    .C(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__o21a_1 _09735_ (.A1(_03930_),
    .A2(_03931_),
    .B1(_03918_),
    .X(_03933_));
 sky130_fd_sc_hd__a211oi_1 _09736_ (.A1(_03789_),
    .A2(_03791_),
    .B1(_03932_),
    .C1(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__a211o_1 _09737_ (.A1(_03789_),
    .A2(_03791_),
    .B1(_03932_),
    .C1(_03933_),
    .X(_03935_));
 sky130_fd_sc_hd__o211ai_1 _09738_ (.A1(_03932_),
    .A2(_03933_),
    .B1(_03789_),
    .C1(_03791_),
    .Y(_03936_));
 sky130_fd_sc_hd__and3_1 _09739_ (.A(_03904_),
    .B(_03935_),
    .C(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__a21oi_1 _09740_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03904_),
    .Y(_03938_));
 sky130_fd_sc_hd__nor3b_2 _09741_ (.A(_03937_),
    .B(_03938_),
    .C_N(_03796_),
    .Y(_03939_));
 sky130_fd_sc_hd__inv_2 _09742_ (.A(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__o21ba_1 _09743_ (.A1(_03937_),
    .A2(_03938_),
    .B1_N(_03796_),
    .X(_03941_));
 sky130_fd_sc_hd__nor4_2 _09744_ (.A(_03893_),
    .B(_03895_),
    .C(_03939_),
    .D(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__or4_2 _09745_ (.A(_03893_),
    .B(_03895_),
    .C(_03939_),
    .D(_03941_),
    .X(_03943_));
 sky130_fd_sc_hd__o22a_1 _09746_ (.A1(_03893_),
    .A2(_03895_),
    .B1(_03939_),
    .B2(_03941_),
    .X(_03944_));
 sky130_fd_sc_hd__a211o_2 _09747_ (.A1(_03798_),
    .A2(_03801_),
    .B1(_03942_),
    .C1(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__o211ai_4 _09748_ (.A1(_03942_),
    .A2(_03944_),
    .B1(_03798_),
    .C1(_03801_),
    .Y(_03946_));
 sky130_fd_sc_hd__o211ai_4 _09749_ (.A1(_03756_),
    .A2(_03758_),
    .B1(_03945_),
    .C1(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__a211o_1 _09750_ (.A1(_03945_),
    .A2(_03946_),
    .B1(_03756_),
    .C1(_03758_),
    .X(_03948_));
 sky130_fd_sc_hd__o211a_1 _09751_ (.A1(_03803_),
    .A2(_03805_),
    .B1(_03947_),
    .C1(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__o211ai_1 _09752_ (.A1(_03803_),
    .A2(_03805_),
    .B1(_03947_),
    .C1(_03948_),
    .Y(_03950_));
 sky130_fd_sc_hd__a211o_1 _09753_ (.A1(_03947_),
    .A2(_03948_),
    .B1(_03803_),
    .C1(_03805_),
    .X(_03951_));
 sky130_fd_sc_hd__and3_1 _09754_ (.A(_03853_),
    .B(_03950_),
    .C(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__a21oi_1 _09755_ (.A1(_03950_),
    .A2(_03951_),
    .B1(_03853_),
    .Y(_03953_));
 sky130_fd_sc_hd__a211oi_2 _09756_ (.A1(_03807_),
    .A2(_03809_),
    .B1(_03952_),
    .C1(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__o211a_1 _09757_ (.A1(_03952_),
    .A2(_03953_),
    .B1(_03807_),
    .C1(_03809_),
    .X(_03955_));
 sky130_fd_sc_hd__nor2_1 _09758_ (.A(_03954_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__and4bb_1 _09759_ (.A_N(_03673_),
    .B_N(_03674_),
    .C(_03811_),
    .D(_03812_),
    .X(_03957_));
 sky130_fd_sc_hd__nand2_1 _09760_ (.A(_03673_),
    .B(_03811_),
    .Y(_03958_));
 sky130_fd_sc_hd__o311a_1 _09761_ (.A1(_03675_),
    .A2(_03676_),
    .A3(_03813_),
    .B1(_03958_),
    .C1(_03812_),
    .X(_03959_));
 sky130_fd_sc_hd__or4b_2 _09762_ (.A(_03323_),
    .B(_03404_),
    .C(_03536_),
    .D_N(_03957_),
    .X(_03960_));
 sky130_fd_sc_hd__nand2_1 _09763_ (.A(_03959_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__or2_1 _09764_ (.A(_03956_),
    .B(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__and2_1 _09765_ (.A(_03956_),
    .B(_03961_),
    .X(_03963_));
 sky130_fd_sc_hd__nand2_1 _09766_ (.A(_03956_),
    .B(_03961_),
    .Y(_03964_));
 sky130_fd_sc_hd__nand3_1 _09767_ (.A(_01869_),
    .B(_01911_),
    .C(_03819_),
    .Y(_03965_));
 sky130_fd_sc_hd__a21o_1 _09768_ (.A1(_01911_),
    .A2(_03819_),
    .B1(_01869_),
    .X(_03966_));
 sky130_fd_sc_hd__a32o_1 _09769_ (.A1(net467),
    .A2(_03965_),
    .A3(_03966_),
    .B1(net485),
    .B2(net3668),
    .X(_03967_));
 sky130_fd_sc_hd__a31o_4 _09770_ (.A1(_02239_),
    .A2(_03962_),
    .A3(_03964_),
    .B1(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__a21oi_4 _09771_ (.A1(net391),
    .A2(_03968_),
    .B1(_03852_),
    .Y(_03969_));
 sky130_fd_sc_hd__nand2_1 _09772_ (.A(net577),
    .B(net3462),
    .Y(_03970_));
 sky130_fd_sc_hd__or2_1 _09773_ (.A(net577),
    .B(net3462),
    .X(_03971_));
 sky130_fd_sc_hd__nand2_1 _09774_ (.A(_03970_),
    .B(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__or3b_1 _09775_ (.A(_01762_),
    .B(_03686_),
    .C_N(_03824_),
    .X(_03973_));
 sky130_fd_sc_hd__o311a_1 _09776_ (.A1(_03687_),
    .A2(_03688_),
    .A3(_03825_),
    .B1(_03973_),
    .C1(_03823_),
    .X(_03974_));
 sky130_fd_sc_hd__o41a_2 _09777_ (.A1(_03418_),
    .A2(_03548_),
    .A3(_03687_),
    .A4(_03825_),
    .B1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__xnor2_1 _09778_ (.A(_03972_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__and2_1 _09779_ (.A(net3537),
    .B(_03697_),
    .X(_03977_));
 sky130_fd_sc_hd__nor2_1 _09780_ (.A(net3537),
    .B(_03697_),
    .Y(_03978_));
 sky130_fd_sc_hd__or3_1 _09781_ (.A(_01958_),
    .B(_03977_),
    .C(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__a21oi_1 _09782_ (.A1(\dpath.btarg_DX.q[20] ),
    .A2(net403),
    .B1(net451),
    .Y(_03980_));
 sky130_fd_sc_hd__o211a_1 _09783_ (.A1(net366),
    .A2(_03976_),
    .B1(_03979_),
    .C1(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__o21ai_1 _09784_ (.A1(net373),
    .A2(_03969_),
    .B1(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__o211a_1 _09785_ (.A1(net3537),
    .A2(net443),
    .B1(_03982_),
    .C1(net844),
    .X(_00656_));
 sky130_fd_sc_hd__mux4_1 _09786_ (.A0(\dpath.RF.R[0][21] ),
    .A1(\dpath.RF.R[1][21] ),
    .A2(\dpath.RF.R[2][21] ),
    .A3(\dpath.RF.R[3][21] ),
    .S0(net568),
    .S1(net549),
    .X(_03983_));
 sky130_fd_sc_hd__mux4_1 _09787_ (.A0(\dpath.RF.R[4][21] ),
    .A1(\dpath.RF.R[5][21] ),
    .A2(\dpath.RF.R[6][21] ),
    .A3(\dpath.RF.R[7][21] ),
    .S0(net568),
    .S1(net549),
    .X(_03984_));
 sky130_fd_sc_hd__o21a_1 _09788_ (.A1(net513),
    .A2(_03984_),
    .B1(net507),
    .X(_03985_));
 sky130_fd_sc_hd__o21ai_1 _09789_ (.A1(net534),
    .A2(_03983_),
    .B1(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__mux4_1 _09790_ (.A0(\dpath.RF.R[12][21] ),
    .A1(\dpath.RF.R[13][21] ),
    .A2(\dpath.RF.R[14][21] ),
    .A3(\dpath.RF.R[15][21] ),
    .S0(net569),
    .S1(net550),
    .X(_03987_));
 sky130_fd_sc_hd__mux4_1 _09791_ (.A0(\dpath.RF.R[8][21] ),
    .A1(\dpath.RF.R[9][21] ),
    .A2(\dpath.RF.R[10][21] ),
    .A3(\dpath.RF.R[11][21] ),
    .S0(net568),
    .S1(net549),
    .X(_03988_));
 sky130_fd_sc_hd__or2_1 _09792_ (.A(net534),
    .B(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__o211a_1 _09793_ (.A1(net513),
    .A2(_03987_),
    .B1(_03989_),
    .C1(net528),
    .X(_03990_));
 sky130_fd_sc_hd__nor2_1 _09794_ (.A(net519),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__mux4_1 _09795_ (.A0(\dpath.RF.R[16][21] ),
    .A1(\dpath.RF.R[17][21] ),
    .A2(\dpath.RF.R[18][21] ),
    .A3(\dpath.RF.R[19][21] ),
    .S0(net568),
    .S1(net549),
    .X(_03992_));
 sky130_fd_sc_hd__nor2_1 _09796_ (.A(net534),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__mux4_1 _09797_ (.A0(\dpath.RF.R[20][21] ),
    .A1(\dpath.RF.R[21][21] ),
    .A2(\dpath.RF.R[22][21] ),
    .A3(\dpath.RF.R[23][21] ),
    .S0(net569),
    .S1(net550),
    .X(_03994_));
 sky130_fd_sc_hd__nor2_1 _09798_ (.A(net513),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__mux4_1 _09799_ (.A0(\dpath.RF.R[28][21] ),
    .A1(\dpath.RF.R[29][21] ),
    .A2(\dpath.RF.R[30][21] ),
    .A3(\dpath.RF.R[31][21] ),
    .S0(net570),
    .S1(net551),
    .X(_03996_));
 sky130_fd_sc_hd__nor2_1 _09800_ (.A(net513),
    .B(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__mux4_1 _09801_ (.A0(\dpath.RF.R[24][21] ),
    .A1(\dpath.RF.R[25][21] ),
    .A2(\dpath.RF.R[26][21] ),
    .A3(\dpath.RF.R[27][21] ),
    .S0(net569),
    .S1(net550),
    .X(_03998_));
 sky130_fd_sc_hd__o21ai_1 _09802_ (.A1(net534),
    .A2(_03998_),
    .B1(net525),
    .Y(_03999_));
 sky130_fd_sc_hd__o32a_1 _09803_ (.A1(net525),
    .A2(_03993_),
    .A3(_03995_),
    .B1(_03997_),
    .B2(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__a221o_1 _09804_ (.A1(_03986_),
    .A2(_03991_),
    .B1(_04000_),
    .B2(net519),
    .C1(net483),
    .X(_04001_));
 sky130_fd_sc_hd__nor2_1 _09805_ (.A(net371),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__mux2_2 _09806_ (.A0(net3658),
    .A1(net14),
    .S(net479),
    .X(_04003_));
 sky130_fd_sc_hd__a221o_1 _09807_ (.A1(net676),
    .A2(net369),
    .B1(net367),
    .B2(_04003_),
    .C1(_04002_),
    .X(_04004_));
 sky130_fd_sc_hd__a22oi_1 _09808_ (.A1(net773),
    .A2(net591),
    .B1(net588),
    .B2(net778),
    .Y(_04005_));
 sky130_fd_sc_hd__and4_1 _09809_ (.A(net778),
    .B(net773),
    .C(net591),
    .D(net588),
    .X(_04006_));
 sky130_fd_sc_hd__o2bb2a_1 _09810_ (.A1_N(net781),
    .A2_N(net586),
    .B1(_04005_),
    .B2(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__and4bb_1 _09811_ (.A_N(_04005_),
    .B_N(_04006_),
    .C(net782),
    .D(net586),
    .X(_04008_));
 sky130_fd_sc_hd__or2_1 _09812_ (.A(_04007_),
    .B(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__nand2_1 _09813_ (.A(_03857_),
    .B(_03859_),
    .Y(_04010_));
 sky130_fd_sc_hd__and2b_1 _09814_ (.A_N(_04009_),
    .B(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__xnor2_1 _09815_ (.A(_04009_),
    .B(_04010_),
    .Y(_04012_));
 sky130_fd_sc_hd__nand2_1 _09816_ (.A(net785),
    .B(net584),
    .Y(_04013_));
 sky130_fd_sc_hd__xor2_1 _09817_ (.A(_04012_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__o21ba_1 _09818_ (.A1(_03855_),
    .A2(_03862_),
    .B1_N(_03861_),
    .X(_04015_));
 sky130_fd_sc_hd__nor2_1 _09819_ (.A(_04014_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__xor2_1 _09820_ (.A(_04014_),
    .B(_04015_),
    .X(_04017_));
 sky130_fd_sc_hd__nand2_1 _09821_ (.A(net789),
    .B(net582),
    .Y(_04018_));
 sky130_fd_sc_hd__xor2_1 _09822_ (.A(_04017_),
    .B(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__a21o_1 _09823_ (.A1(_03909_),
    .A2(_03916_),
    .B1(_03915_),
    .X(_04020_));
 sky130_fd_sc_hd__nand2_1 _09824_ (.A(_03874_),
    .B(_03876_),
    .Y(_04021_));
 sky130_fd_sc_hd__a22o_1 _09825_ (.A1(net761),
    .A2(net599),
    .B1(net595),
    .B2(net766),
    .X(_04022_));
 sky130_fd_sc_hd__nand4_1 _09826_ (.A(net766),
    .B(net761),
    .C(net599),
    .D(net595),
    .Y(_04023_));
 sky130_fd_sc_hd__a22oi_2 _09827_ (.A1(net769),
    .A2(net593),
    .B1(_04022_),
    .B2(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__and4_1 _09828_ (.A(net769),
    .B(net593),
    .C(_04022_),
    .D(_04023_),
    .X(_04025_));
 sky130_fd_sc_hd__a211o_2 _09829_ (.A1(_03906_),
    .A2(_03907_),
    .B1(_04024_),
    .C1(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__o211ai_2 _09830_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_03906_),
    .C1(_03907_),
    .Y(_04027_));
 sky130_fd_sc_hd__nand3_2 _09831_ (.A(_04021_),
    .B(_04026_),
    .C(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__a21o_1 _09832_ (.A1(_04026_),
    .A2(_04027_),
    .B1(_04021_),
    .X(_04029_));
 sky130_fd_sc_hd__and3_2 _09833_ (.A(_04020_),
    .B(_04028_),
    .C(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__a21oi_2 _09834_ (.A1(_04028_),
    .A2(_04029_),
    .B1(_04020_),
    .Y(_04031_));
 sky130_fd_sc_hd__a211oi_4 _09835_ (.A1(_03877_),
    .A2(_03879_),
    .B1(_04030_),
    .C1(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__o211a_1 _09836_ (.A1(_04030_),
    .A2(_04031_),
    .B1(_03877_),
    .C1(_03879_),
    .X(_04033_));
 sky130_fd_sc_hd__a211oi_2 _09837_ (.A1(_03882_),
    .A2(_03884_),
    .B1(_04032_),
    .C1(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__o211a_1 _09838_ (.A1(_04032_),
    .A2(_04033_),
    .B1(_03882_),
    .C1(_03884_),
    .X(_04035_));
 sky130_fd_sc_hd__or3_1 _09839_ (.A(_04019_),
    .B(_04034_),
    .C(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__o21ai_1 _09840_ (.A1(_04034_),
    .A2(_04035_),
    .B1(_04019_),
    .Y(_04037_));
 sky130_fd_sc_hd__and3_2 _09841_ (.A(_03934_),
    .B(_04036_),
    .C(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__a21oi_2 _09842_ (.A1(_04036_),
    .A2(_04037_),
    .B1(_03934_),
    .Y(_04039_));
 sky130_fd_sc_hd__a211oi_4 _09843_ (.A1(_03886_),
    .A2(_03888_),
    .B1(_04038_),
    .C1(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__o211a_1 _09844_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_03886_),
    .C1(_03888_),
    .X(_04041_));
 sky130_fd_sc_hd__a22oi_1 _09845_ (.A1(net649),
    .A2(\dpath.alu.adder.in1[20] ),
    .B1(net724),
    .B2(net653),
    .Y(_04042_));
 sky130_fd_sc_hd__and4_1 _09846_ (.A(net653),
    .B(net649),
    .C(net725),
    .D(net724),
    .X(_04043_));
 sky130_fd_sc_hd__or2_1 _09847_ (.A(_04042_),
    .B(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__and2_1 _09848_ (.A(net635),
    .B(net731),
    .X(_04045_));
 sky130_fd_sc_hd__a22o_1 _09849_ (.A1(net639),
    .A2(net729),
    .B1(net727),
    .B2(net645),
    .X(_04046_));
 sky130_fd_sc_hd__nand4_1 _09850_ (.A(net645),
    .B(net639),
    .C(net729),
    .D(net727),
    .Y(_04047_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(_04046_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__xnor2_2 _09852_ (.A(_04045_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__nand2b_1 _09853_ (.A_N(_04044_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__xnor2_2 _09854_ (.A(_04044_),
    .B(_04049_),
    .Y(_04051_));
 sky130_fd_sc_hd__nand2b_1 _09855_ (.A_N(_03903_),
    .B(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__xnor2_1 _09856_ (.A(_03903_),
    .B(_04051_),
    .Y(_04053_));
 sky130_fd_sc_hd__a22o_1 _09857_ (.A1(net751),
    .A2(net608),
    .B1(net606),
    .B2(net754),
    .X(_04054_));
 sky130_fd_sc_hd__and3_1 _09858_ (.A(net754),
    .B(net751),
    .C(net608),
    .X(_04055_));
 sky130_fd_sc_hd__a21bo_1 _09859_ (.A1(net606),
    .A2(_04055_),
    .B1_N(_04054_),
    .X(_04056_));
 sky130_fd_sc_hd__nand2_2 _09860_ (.A(net757),
    .B(net603),
    .Y(_04057_));
 sky130_fd_sc_hd__xnor2_4 _09861_ (.A(_04056_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__a22o_1 _09862_ (.A1(net613),
    .A2(net744),
    .B1(net740),
    .B2(net616),
    .X(_04059_));
 sky130_fd_sc_hd__and4_1 _09863_ (.A(net616),
    .B(net615),
    .C(net746),
    .D(net742),
    .X(_04060_));
 sky130_fd_sc_hd__nand4_2 _09864_ (.A(net616),
    .B(net615),
    .C(net744),
    .D(net740),
    .Y(_04061_));
 sky130_fd_sc_hd__and4_1 _09865_ (.A(net611),
    .B(net750),
    .C(_04059_),
    .D(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__nand4_1 _09866_ (.A(net611),
    .B(net748),
    .C(_04059_),
    .D(_04061_),
    .Y(_04063_));
 sky130_fd_sc_hd__a22o_1 _09867_ (.A1(net611),
    .A2(net748),
    .B1(_04059_),
    .B2(_04061_),
    .X(_04064_));
 sky130_fd_sc_hd__a21bo_1 _09868_ (.A1(_03910_),
    .A2(_03911_),
    .B1_N(_03912_),
    .X(_04065_));
 sky130_fd_sc_hd__and3_1 _09869_ (.A(_04063_),
    .B(_04064_),
    .C(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__a21oi_1 _09870_ (.A1(_04063_),
    .A2(_04064_),
    .B1(_04065_),
    .Y(_04067_));
 sky130_fd_sc_hd__nor2_2 _09871_ (.A(_04066_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__xnor2_4 _09872_ (.A(_04058_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__a41o_1 _09873_ (.A1(net635),
    .A2(net631),
    .A3(net734),
    .A4(net732),
    .B1(_03924_),
    .X(_04070_));
 sky130_fd_sc_hd__a31o_1 _09874_ (.A1(net639),
    .A2(net731),
    .A3(_03897_),
    .B1(_03899_),
    .X(_04071_));
 sky130_fd_sc_hd__a22o_1 _09875_ (.A1(net627),
    .A2(net734),
    .B1(net732),
    .B2(net631),
    .X(_04072_));
 sky130_fd_sc_hd__nand4_2 _09876_ (.A(net631),
    .B(net627),
    .C(\dpath.alu.adder.in1[15] ),
    .D(\dpath.alu.adder.in1[16] ),
    .Y(_04073_));
 sky130_fd_sc_hd__a22o_1 _09877_ (.A1(net623),
    .A2(net737),
    .B1(_04072_),
    .B2(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__nand4_2 _09878_ (.A(net623),
    .B(net737),
    .C(_04072_),
    .D(_04073_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand3_1 _09879_ (.A(_04071_),
    .B(_04074_),
    .C(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__a21o_1 _09880_ (.A1(_04074_),
    .A2(_04075_),
    .B1(_04071_),
    .X(_04077_));
 sky130_fd_sc_hd__and3_1 _09881_ (.A(_04070_),
    .B(_04076_),
    .C(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__a21oi_1 _09882_ (.A1(_04076_),
    .A2(_04077_),
    .B1(_04070_),
    .Y(_04079_));
 sky130_fd_sc_hd__or2_1 _09883_ (.A(_04078_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__a21o_1 _09884_ (.A1(_03926_),
    .A2(_03928_),
    .B1(_04080_),
    .X(_04081_));
 sky130_fd_sc_hd__inv_2 _09885_ (.A(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand3_2 _09886_ (.A(_03926_),
    .B(_03928_),
    .C(_04080_),
    .Y(_04083_));
 sky130_fd_sc_hd__and3_1 _09887_ (.A(_04069_),
    .B(_04081_),
    .C(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__nand3_2 _09888_ (.A(_04069_),
    .B(_04081_),
    .C(_04083_),
    .Y(_04085_));
 sky130_fd_sc_hd__a21o_1 _09889_ (.A1(_04081_),
    .A2(_04083_),
    .B1(_04069_),
    .X(_04086_));
 sky130_fd_sc_hd__o211ai_4 _09890_ (.A1(_03930_),
    .A2(_03932_),
    .B1(_04085_),
    .C1(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__a211o_1 _09891_ (.A1(_04085_),
    .A2(_04086_),
    .B1(_03930_),
    .C1(_03932_),
    .X(_04088_));
 sky130_fd_sc_hd__and3_2 _09892_ (.A(_04053_),
    .B(_04087_),
    .C(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__a21oi_2 _09893_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_04053_),
    .Y(_04090_));
 sky130_fd_sc_hd__nor3b_4 _09894_ (.A(_04089_),
    .B(_04090_),
    .C_N(_03937_),
    .Y(_04091_));
 sky130_fd_sc_hd__o21ba_1 _09895_ (.A1(_04089_),
    .A2(_04090_),
    .B1_N(_03937_),
    .X(_04092_));
 sky130_fd_sc_hd__nor4_4 _09896_ (.A(_04040_),
    .B(_04041_),
    .C(_04091_),
    .D(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__o22a_1 _09897_ (.A1(_04040_),
    .A2(_04041_),
    .B1(_04091_),
    .B2(_04092_),
    .X(_04094_));
 sky130_fd_sc_hd__a211oi_4 _09898_ (.A1(_03940_),
    .A2(_03943_),
    .B1(_04093_),
    .C1(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__o211a_1 _09899_ (.A1(_04093_),
    .A2(_04094_),
    .B1(_03940_),
    .C1(_03943_),
    .X(_04096_));
 sky130_fd_sc_hd__a211oi_4 _09900_ (.A1(_03891_),
    .A2(_03894_),
    .B1(_04095_),
    .C1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__o211a_1 _09901_ (.A1(_04095_),
    .A2(_04096_),
    .B1(_03891_),
    .C1(_03894_),
    .X(_04098_));
 sky130_fd_sc_hd__a211oi_4 _09902_ (.A1(_03945_),
    .A2(_03947_),
    .B1(_04097_),
    .C1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__inv_2 _09903_ (.A(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__o211a_1 _09904_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_03945_),
    .C1(_03947_),
    .X(_04101_));
 sky130_fd_sc_hd__a211o_2 _09905_ (.A1(_03865_),
    .A2(_03868_),
    .B1(_04099_),
    .C1(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__o211ai_2 _09906_ (.A1(_04099_),
    .A2(_04101_),
    .B1(_03865_),
    .C1(_03868_),
    .Y(_04103_));
 sky130_fd_sc_hd__o211a_1 _09907_ (.A1(_03949_),
    .A2(_03952_),
    .B1(_04102_),
    .C1(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__a211oi_2 _09908_ (.A1(_04102_),
    .A2(_04103_),
    .B1(_03949_),
    .C1(_03952_),
    .Y(_04105_));
 sky130_fd_sc_hd__nor2_1 _09909_ (.A(_04104_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__nor2_1 _09910_ (.A(_03954_),
    .B(_03963_),
    .Y(_04107_));
 sky130_fd_sc_hd__xnor2_1 _09911_ (.A(_04106_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__or2_1 _09912_ (.A(net3686),
    .B(_02071_),
    .X(_04109_));
 sky130_fd_sc_hd__o211a_1 _09913_ (.A1(net486),
    .A2(_04108_),
    .B1(_04109_),
    .C1(net468),
    .X(_04110_));
 sky130_fd_sc_hd__nand3_1 _09914_ (.A(_01867_),
    .B(_01881_),
    .C(_03966_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21o_1 _09915_ (.A1(_01867_),
    .A2(_03966_),
    .B1(_01881_),
    .X(_04112_));
 sky130_fd_sc_hd__a31o_4 _09916_ (.A1(_02101_),
    .A2(_04111_),
    .A3(_04112_),
    .B1(_04110_),
    .X(_04113_));
 sky130_fd_sc_hd__a21oi_4 _09917_ (.A1(net391),
    .A2(_04113_),
    .B1(_04004_),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _09918_ (.A(net373),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__xor2_1 _09919_ (.A(net577),
    .B(net3455),
    .X(_04116_));
 sky130_fd_sc_hd__o21ai_1 _09920_ (.A1(_03972_),
    .A2(_03975_),
    .B1(_03970_),
    .Y(_04117_));
 sky130_fd_sc_hd__xnor2_1 _09921_ (.A(_04116_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__nor2_1 _09922_ (.A(net366),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _09923_ (.A(net241),
    .B(_03977_),
    .Y(_04120_));
 sky130_fd_sc_hd__o211a_1 _09924_ (.A1(net241),
    .A2(_03977_),
    .B1(_04120_),
    .C1(net362),
    .X(_04121_));
 sky130_fd_sc_hd__a2111o_1 _09925_ (.A1(net3372),
    .A2(net403),
    .B1(net451),
    .C1(_04119_),
    .D1(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__o221a_1 _09926_ (.A1(net241),
    .A2(net443),
    .B1(_04115_),
    .B2(net3373),
    .C1(net844),
    .X(_00657_));
 sky130_fd_sc_hd__xnor2_1 _09927_ (.A(net577),
    .B(net3466),
    .Y(_04123_));
 sky130_fd_sc_hd__o21ai_1 _09928_ (.A1(net3455),
    .A2(net3462),
    .B1(net577),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2b_1 _09929_ (.A_N(_03972_),
    .B(_04116_),
    .Y(_04125_));
 sky130_fd_sc_hd__or2_1 _09930_ (.A(_03975_),
    .B(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__a21oi_1 _09931_ (.A1(_04124_),
    .A2(_04126_),
    .B1(_04123_),
    .Y(_04127_));
 sky130_fd_sc_hd__and3_1 _09932_ (.A(_04123_),
    .B(_04124_),
    .C(_04126_),
    .X(_04128_));
 sky130_fd_sc_hd__or2_1 _09933_ (.A(_04127_),
    .B(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__nor2_1 _09934_ (.A(net366),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__mux4_1 _09935_ (.A0(\dpath.RF.R[0][22] ),
    .A1(\dpath.RF.R[1][22] ),
    .A2(\dpath.RF.R[2][22] ),
    .A3(\dpath.RF.R[3][22] ),
    .S0(net571),
    .S1(net552),
    .X(_04131_));
 sky130_fd_sc_hd__mux4_1 _09936_ (.A0(\dpath.RF.R[4][22] ),
    .A1(\dpath.RF.R[5][22] ),
    .A2(\dpath.RF.R[6][22] ),
    .A3(\dpath.RF.R[7][22] ),
    .S0(net571),
    .S1(net552),
    .X(_04132_));
 sky130_fd_sc_hd__o21a_1 _09937_ (.A1(net516),
    .A2(_04132_),
    .B1(net506),
    .X(_04133_));
 sky130_fd_sc_hd__o21ai_1 _09938_ (.A1(net537),
    .A2(_04131_),
    .B1(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__mux4_1 _09939_ (.A0(\dpath.RF.R[12][22] ),
    .A1(\dpath.RF.R[13][22] ),
    .A2(\dpath.RF.R[14][22] ),
    .A3(\dpath.RF.R[15][22] ),
    .S0(net571),
    .S1(net552),
    .X(_04135_));
 sky130_fd_sc_hd__mux4_1 _09940_ (.A0(\dpath.RF.R[8][22] ),
    .A1(\dpath.RF.R[9][22] ),
    .A2(\dpath.RF.R[10][22] ),
    .A3(\dpath.RF.R[11][22] ),
    .S0(net567),
    .S1(net548),
    .X(_04136_));
 sky130_fd_sc_hd__or2_1 _09941_ (.A(net535),
    .B(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__o211a_1 _09942_ (.A1(net514),
    .A2(_04135_),
    .B1(_04137_),
    .C1(net527),
    .X(_04138_));
 sky130_fd_sc_hd__nor2_1 _09943_ (.A(net520),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__mux4_1 _09944_ (.A0(\dpath.RF.R[16][22] ),
    .A1(\dpath.RF.R[17][22] ),
    .A2(\dpath.RF.R[18][22] ),
    .A3(\dpath.RF.R[19][22] ),
    .S0(net571),
    .S1(net552),
    .X(_04140_));
 sky130_fd_sc_hd__nor2_1 _09945_ (.A(net537),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__mux4_1 _09946_ (.A0(\dpath.RF.R[20][22] ),
    .A1(\dpath.RF.R[21][22] ),
    .A2(\dpath.RF.R[22][22] ),
    .A3(\dpath.RF.R[23][22] ),
    .S0(net571),
    .S1(net552),
    .X(_04142_));
 sky130_fd_sc_hd__nor2_1 _09947_ (.A(net516),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__mux4_1 _09948_ (.A0(\dpath.RF.R[28][22] ),
    .A1(\dpath.RF.R[29][22] ),
    .A2(\dpath.RF.R[30][22] ),
    .A3(\dpath.RF.R[31][22] ),
    .S0(net572),
    .S1(net553),
    .X(_04144_));
 sky130_fd_sc_hd__nor2_1 _09949_ (.A(net516),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__mux4_1 _09950_ (.A0(\dpath.RF.R[24][22] ),
    .A1(\dpath.RF.R[25][22] ),
    .A2(\dpath.RF.R[26][22] ),
    .A3(\dpath.RF.R[27][22] ),
    .S0(net572),
    .S1(net553),
    .X(_04146_));
 sky130_fd_sc_hd__o21ai_1 _09951_ (.A1(net537),
    .A2(_04146_),
    .B1(net527),
    .Y(_04147_));
 sky130_fd_sc_hd__o32a_1 _09952_ (.A1(net527),
    .A2(_04141_),
    .A3(_04143_),
    .B1(_04145_),
    .B2(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__a221o_1 _09953_ (.A1(_04134_),
    .A2(_04139_),
    .B1(_04148_),
    .B2(net520),
    .C1(net483),
    .X(_04149_));
 sky130_fd_sc_hd__nor2_1 _09954_ (.A(net371),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__mux2_2 _09955_ (.A0(net3622),
    .A1(net15),
    .S(net479),
    .X(_04151_));
 sky130_fd_sc_hd__a221o_1 _09956_ (.A1(net673),
    .A2(net369),
    .B1(net367),
    .B2(_04151_),
    .C1(_04150_),
    .X(_04152_));
 sky130_fd_sc_hd__a31o_1 _09957_ (.A1(net789),
    .A2(net582),
    .A3(_04017_),
    .B1(_04016_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2b_1 _09958_ (.A_N(_04034_),
    .B(_04036_),
    .Y(_04154_));
 sky130_fd_sc_hd__a22oi_1 _09959_ (.A1(net773),
    .A2(net588),
    .B1(net586),
    .B2(net778),
    .Y(_04155_));
 sky130_fd_sc_hd__and4_1 _09960_ (.A(net778),
    .B(net773),
    .C(net588),
    .D(net586),
    .X(_04156_));
 sky130_fd_sc_hd__o2bb2a_1 _09961_ (.A1_N(net782),
    .A2_N(net584),
    .B1(_04155_),
    .B2(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__and4bb_1 _09962_ (.A_N(_04155_),
    .B_N(_04156_),
    .C(net782),
    .D(net584),
    .X(_04158_));
 sky130_fd_sc_hd__or2_1 _09963_ (.A(_04157_),
    .B(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__or2_1 _09964_ (.A(_04006_),
    .B(_04008_),
    .X(_04160_));
 sky130_fd_sc_hd__and2b_1 _09965_ (.A_N(_04159_),
    .B(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__xnor2_2 _09966_ (.A(_04159_),
    .B(_04160_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(\dpath.alu.adder.in1[1] ),
    .B(net582),
    .Y(_04163_));
 sky130_fd_sc_hd__xnor2_2 _09968_ (.A(_04162_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__a31o_1 _09969_ (.A1(\dpath.alu.adder.in1[1] ),
    .A2(net584),
    .A3(_04012_),
    .B1(_04011_),
    .X(_04165_));
 sky130_fd_sc_hd__nand2_1 _09970_ (.A(_04164_),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__xor2_2 _09971_ (.A(_04164_),
    .B(_04165_),
    .X(_04167_));
 sky130_fd_sc_hd__nand2_1 _09972_ (.A(\dpath.alu.adder.in1[0] ),
    .B(net580),
    .Y(_04168_));
 sky130_fd_sc_hd__nand3_2 _09973_ (.A(net789),
    .B(net580),
    .C(_04167_),
    .Y(_04169_));
 sky130_fd_sc_hd__xor2_1 _09974_ (.A(_04167_),
    .B(_04168_),
    .X(_04170_));
 sky130_fd_sc_hd__o21bai_2 _09975_ (.A1(_04058_),
    .A2(_04067_),
    .B1_N(_04066_),
    .Y(_04171_));
 sky130_fd_sc_hd__a41o_1 _09976_ (.A1(net766),
    .A2(net761),
    .A3(net600),
    .A4(net597),
    .B1(_04025_),
    .X(_04172_));
 sky130_fd_sc_hd__a32o_1 _09977_ (.A1(net757),
    .A2(net603),
    .A3(_04054_),
    .B1(_04055_),
    .B2(net606),
    .X(_04173_));
 sky130_fd_sc_hd__a22o_1 _09978_ (.A1(net761),
    .A2(net597),
    .B1(net594),
    .B2(net766),
    .X(_04174_));
 sky130_fd_sc_hd__nand4_2 _09979_ (.A(net766),
    .B(net761),
    .C(net597),
    .D(net594),
    .Y(_04175_));
 sky130_fd_sc_hd__a22o_1 _09980_ (.A1(net769),
    .A2(net589),
    .B1(_04174_),
    .B2(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__nand4_2 _09981_ (.A(net769),
    .B(net589),
    .C(_04174_),
    .D(_04175_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand3_4 _09982_ (.A(_04173_),
    .B(_04176_),
    .C(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__a21o_1 _09983_ (.A1(_04176_),
    .A2(_04177_),
    .B1(_04173_),
    .X(_04179_));
 sky130_fd_sc_hd__nand3_4 _09984_ (.A(_04172_),
    .B(_04178_),
    .C(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__a21o_1 _09985_ (.A1(_04178_),
    .A2(_04179_),
    .B1(_04172_),
    .X(_04181_));
 sky130_fd_sc_hd__and3_1 _09986_ (.A(_04171_),
    .B(_04180_),
    .C(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__nand3_2 _09987_ (.A(_04171_),
    .B(_04180_),
    .C(_04181_),
    .Y(_04183_));
 sky130_fd_sc_hd__a21oi_1 _09988_ (.A1(_04180_),
    .A2(_04181_),
    .B1(_04171_),
    .Y(_04184_));
 sky130_fd_sc_hd__a211o_2 _09989_ (.A1(_04026_),
    .A2(_04028_),
    .B1(_04182_),
    .C1(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__o211ai_2 _09990_ (.A1(_04182_),
    .A2(_04184_),
    .B1(_04026_),
    .C1(_04028_),
    .Y(_04186_));
 sky130_fd_sc_hd__o211a_2 _09991_ (.A1(_04030_),
    .A2(_04032_),
    .B1(_04185_),
    .C1(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__a211oi_2 _09992_ (.A1(_04185_),
    .A2(_04186_),
    .B1(_04030_),
    .C1(_04032_),
    .Y(_04188_));
 sky130_fd_sc_hd__nor3_2 _09993_ (.A(_04170_),
    .B(_04187_),
    .C(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__o21a_1 _09994_ (.A1(_04187_),
    .A2(_04188_),
    .B1(_04170_),
    .X(_04190_));
 sky130_fd_sc_hd__or3_2 _09995_ (.A(_04087_),
    .B(_04189_),
    .C(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__o21ai_1 _09996_ (.A1(_04189_),
    .A2(_04190_),
    .B1(_04087_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand3_2 _09997_ (.A(_04154_),
    .B(_04191_),
    .C(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__a21o_1 _09998_ (.A1(_04191_),
    .A2(_04192_),
    .B1(_04154_),
    .X(_04194_));
 sky130_fd_sc_hd__a22oi_1 _09999_ (.A1(net648),
    .A2(net724),
    .B1(\dpath.alu.adder.in1[22] ),
    .B2(net653),
    .Y(_04195_));
 sky130_fd_sc_hd__and4_1 _10000_ (.A(net653),
    .B(net648),
    .C(net724),
    .D(\dpath.alu.adder.in1[22] ),
    .X(_04196_));
 sky130_fd_sc_hd__o2bb2a_1 _10001_ (.A1_N(net645),
    .A2_N(\dpath.alu.adder.in1[20] ),
    .B1(_04195_),
    .B2(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__and4bb_1 _10002_ (.A_N(_04195_),
    .B_N(_04196_),
    .C(net645),
    .D(\dpath.alu.adder.in1[20] ),
    .X(_04198_));
 sky130_fd_sc_hd__nor2_1 _10003_ (.A(_04197_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__and2_1 _10004_ (.A(_04043_),
    .B(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__xnor2_2 _10005_ (.A(_04043_),
    .B(_04199_),
    .Y(_04201_));
 sky130_fd_sc_hd__a22o_1 _10006_ (.A1(net635),
    .A2(net729),
    .B1(net727),
    .B2(net639),
    .X(_04202_));
 sky130_fd_sc_hd__and4_1 _10007_ (.A(net639),
    .B(net635),
    .C(net729),
    .D(net727),
    .X(_04203_));
 sky130_fd_sc_hd__nand4_1 _10008_ (.A(\dpath.alu.adder.in0[3] ),
    .B(net635),
    .C(net729),
    .D(net727),
    .Y(_04204_));
 sky130_fd_sc_hd__a22oi_1 _10009_ (.A1(net631),
    .A2(net731),
    .B1(_04202_),
    .B2(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__and4_1 _10010_ (.A(net631),
    .B(net731),
    .C(_04202_),
    .D(_04204_),
    .X(_04206_));
 sky130_fd_sc_hd__or2_1 _10011_ (.A(_04205_),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(_04201_),
    .B(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__xor2_2 _10013_ (.A(_04201_),
    .B(_04207_),
    .X(_04209_));
 sky130_fd_sc_hd__nand2b_1 _10014_ (.A_N(_04050_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_2 _10015_ (.A(_04050_),
    .B(_04209_),
    .Y(_04211_));
 sky130_fd_sc_hd__a22o_1 _10016_ (.A1(net752),
    .A2(net604),
    .B1(net601),
    .B2(net755),
    .X(_04212_));
 sky130_fd_sc_hd__nand4_4 _10017_ (.A(net755),
    .B(net752),
    .C(net604),
    .D(net601),
    .Y(_04213_));
 sky130_fd_sc_hd__a22o_1 _10018_ (.A1(net758),
    .A2(net598),
    .B1(_04212_),
    .B2(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__nand4_2 _10019_ (.A(net758),
    .B(net598),
    .C(_04212_),
    .D(_04213_),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_1 _10020_ (.A(_04214_),
    .B(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__a22oi_2 _10021_ (.A1(net611),
    .A2(net746),
    .B1(net742),
    .B2(net615),
    .Y(_04217_));
 sky130_fd_sc_hd__and4_1 _10022_ (.A(net615),
    .B(net611),
    .C(net746),
    .D(net742),
    .X(_04218_));
 sky130_fd_sc_hd__nor3_1 _10023_ (.A(_01885_),
    .B(_04217_),
    .C(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__or3_1 _10024_ (.A(_01885_),
    .B(_04217_),
    .C(_04218_),
    .X(_04220_));
 sky130_fd_sc_hd__o21ai_1 _10025_ (.A1(_04217_),
    .A2(_04218_),
    .B1(_01885_),
    .Y(_04221_));
 sky130_fd_sc_hd__o211a_1 _10026_ (.A1(_04060_),
    .A2(_04062_),
    .B1(_04220_),
    .C1(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__a211o_1 _10027_ (.A1(_04220_),
    .A2(_04221_),
    .B1(_04060_),
    .C1(_04062_),
    .X(_04223_));
 sky130_fd_sc_hd__and2b_1 _10028_ (.A_N(_04222_),
    .B(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__xnor2_2 _10029_ (.A(_04216_),
    .B(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__nand2_1 _10030_ (.A(_04073_),
    .B(_04075_),
    .Y(_04226_));
 sky130_fd_sc_hd__a21bo_1 _10031_ (.A1(_04045_),
    .A2(_04046_),
    .B1_N(_04047_),
    .X(_04227_));
 sky130_fd_sc_hd__a22o_1 _10032_ (.A1(net622),
    .A2(\dpath.alu.adder.in1[15] ),
    .B1(\dpath.alu.adder.in1[16] ),
    .B2(net627),
    .X(_04228_));
 sky130_fd_sc_hd__nand4_1 _10033_ (.A(net627),
    .B(net623),
    .C(net735),
    .D(net733),
    .Y(_04229_));
 sky130_fd_sc_hd__a22o_1 _10034_ (.A1(net619),
    .A2(net737),
    .B1(_04228_),
    .B2(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__nand4_1 _10035_ (.A(net619),
    .B(net737),
    .C(_04228_),
    .D(_04229_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand3_1 _10036_ (.A(_04227_),
    .B(_04230_),
    .C(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__a21o_1 _10037_ (.A1(_04230_),
    .A2(_04231_),
    .B1(_04227_),
    .X(_04233_));
 sky130_fd_sc_hd__nand3_1 _10038_ (.A(_04226_),
    .B(_04232_),
    .C(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__a21o_1 _10039_ (.A1(_04232_),
    .A2(_04233_),
    .B1(_04226_),
    .X(_04235_));
 sky130_fd_sc_hd__a21bo_1 _10040_ (.A1(_04070_),
    .A2(_04077_),
    .B1_N(_04076_),
    .X(_04236_));
 sky130_fd_sc_hd__and3_1 _10041_ (.A(_04234_),
    .B(_04235_),
    .C(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__nand3_1 _10042_ (.A(_04234_),
    .B(_04235_),
    .C(_04236_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21o_1 _10043_ (.A1(_04234_),
    .A2(_04235_),
    .B1(_04236_),
    .X(_04239_));
 sky130_fd_sc_hd__and3_2 _10044_ (.A(_04225_),
    .B(_04238_),
    .C(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__a21oi_1 _10045_ (.A1(_04238_),
    .A2(_04239_),
    .B1(_04225_),
    .Y(_04241_));
 sky130_fd_sc_hd__or3_4 _10046_ (.A(_04052_),
    .B(_04240_),
    .C(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__o21ai_2 _10047_ (.A1(_04240_),
    .A2(_04241_),
    .B1(_04052_),
    .Y(_04243_));
 sky130_fd_sc_hd__o211ai_4 _10048_ (.A1(_04082_),
    .A2(_04084_),
    .B1(_04242_),
    .C1(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__a211o_1 _10049_ (.A1(_04242_),
    .A2(_04243_),
    .B1(_04082_),
    .C1(_04084_),
    .X(_04245_));
 sky130_fd_sc_hd__nand3_2 _10050_ (.A(_04211_),
    .B(_04244_),
    .C(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__a21o_1 _10051_ (.A1(_04244_),
    .A2(_04245_),
    .B1(_04211_),
    .X(_04247_));
 sky130_fd_sc_hd__nand3_2 _10052_ (.A(_04089_),
    .B(_04246_),
    .C(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__inv_2 _10053_ (.A(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__a21o_1 _10054_ (.A1(_04246_),
    .A2(_04247_),
    .B1(_04089_),
    .X(_04250_));
 sky130_fd_sc_hd__and4_1 _10055_ (.A(_04193_),
    .B(_04194_),
    .C(_04248_),
    .D(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__nand4_2 _10056_ (.A(_04193_),
    .B(_04194_),
    .C(_04248_),
    .D(_04250_),
    .Y(_04252_));
 sky130_fd_sc_hd__a22o_1 _10057_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04248_),
    .B2(_04250_),
    .X(_04253_));
 sky130_fd_sc_hd__o211ai_4 _10058_ (.A1(_04091_),
    .A2(_04093_),
    .B1(_04252_),
    .C1(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__a211o_1 _10059_ (.A1(_04252_),
    .A2(_04253_),
    .B1(_04091_),
    .C1(_04093_),
    .X(_04255_));
 sky130_fd_sc_hd__o211ai_4 _10060_ (.A1(_04038_),
    .A2(_04040_),
    .B1(_04254_),
    .C1(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__a211o_1 _10061_ (.A1(_04254_),
    .A2(_04255_),
    .B1(_04038_),
    .C1(_04040_),
    .X(_04257_));
 sky130_fd_sc_hd__o211ai_4 _10062_ (.A1(_04095_),
    .A2(_04097_),
    .B1(_04256_),
    .C1(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__a211o_1 _10063_ (.A1(_04256_),
    .A2(_04257_),
    .B1(_04095_),
    .C1(_04097_),
    .X(_04259_));
 sky130_fd_sc_hd__and3_1 _10064_ (.A(_04153_),
    .B(_04258_),
    .C(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__nand3_1 _10065_ (.A(_04153_),
    .B(_04258_),
    .C(_04259_),
    .Y(_04261_));
 sky130_fd_sc_hd__a21oi_1 _10066_ (.A1(_04258_),
    .A2(_04259_),
    .B1(_04153_),
    .Y(_04262_));
 sky130_fd_sc_hd__a211oi_2 _10067_ (.A1(_04100_),
    .A2(_04102_),
    .B1(_04260_),
    .C1(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__o211a_1 _10068_ (.A1(_04260_),
    .A2(_04262_),
    .B1(_04100_),
    .C1(_04102_),
    .X(_04264_));
 sky130_fd_sc_hd__or2_1 _10069_ (.A(_04263_),
    .B(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__o21bai_1 _10070_ (.A1(_03954_),
    .A2(_04104_),
    .B1_N(_04105_),
    .Y(_04266_));
 sky130_fd_sc_hd__or3b_1 _10071_ (.A(_04104_),
    .B(_04105_),
    .C_N(_03956_),
    .X(_04267_));
 sky130_fd_sc_hd__a21o_1 _10072_ (.A1(_03959_),
    .A2(_03960_),
    .B1(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__and3_1 _10073_ (.A(_04265_),
    .B(_04266_),
    .C(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__a21oi_1 _10074_ (.A1(_04266_),
    .A2(_04268_),
    .B1(_04265_),
    .Y(_04270_));
 sky130_fd_sc_hd__or3_2 _10075_ (.A(_02240_),
    .B(_04269_),
    .C(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__a21o_1 _10076_ (.A1(_01879_),
    .A2(_04112_),
    .B1(_01922_),
    .X(_04272_));
 sky130_fd_sc_hd__nand2_1 _10077_ (.A(net467),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a31o_1 _10078_ (.A1(_01879_),
    .A2(_01922_),
    .A3(_04112_),
    .B1(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__o211ai_4 _10079_ (.A1(_01786_),
    .A2(net484),
    .B1(_04271_),
    .C1(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__a21oi_4 _10080_ (.A1(net391),
    .A2(_04275_),
    .B1(_04152_),
    .Y(_04276_));
 sky130_fd_sc_hd__nor2_1 _10081_ (.A(net374),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _10082_ (.A(_01761_),
    .B(_04120_),
    .Y(_04278_));
 sky130_fd_sc_hd__a211oi_1 _10083_ (.A1(_01761_),
    .A2(_04120_),
    .B1(_04278_),
    .C1(_01958_),
    .Y(_04279_));
 sky130_fd_sc_hd__a2111o_1 _10084_ (.A1(net3396),
    .A2(net404),
    .B1(net451),
    .C1(_04130_),
    .D1(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__o221a_1 _10085_ (.A1(net242),
    .A2(net443),
    .B1(_04277_),
    .B2(net3397),
    .C1(net851),
    .X(_00658_));
 sky130_fd_sc_hd__mux4_1 _10086_ (.A0(\dpath.RF.R[0][23] ),
    .A1(\dpath.RF.R[1][23] ),
    .A2(\dpath.RF.R[2][23] ),
    .A3(\dpath.RF.R[3][23] ),
    .S0(net567),
    .S1(net548),
    .X(_04281_));
 sky130_fd_sc_hd__mux4_1 _10087_ (.A0(\dpath.RF.R[4][23] ),
    .A1(\dpath.RF.R[5][23] ),
    .A2(\dpath.RF.R[6][23] ),
    .A3(\dpath.RF.R[7][23] ),
    .S0(net567),
    .S1(net548),
    .X(_04282_));
 sky130_fd_sc_hd__o21a_1 _10088_ (.A1(net513),
    .A2(_04282_),
    .B1(net507),
    .X(_04283_));
 sky130_fd_sc_hd__o21ai_1 _10089_ (.A1(net535),
    .A2(_04281_),
    .B1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__mux4_1 _10090_ (.A0(\dpath.RF.R[12][23] ),
    .A1(\dpath.RF.R[13][23] ),
    .A2(\dpath.RF.R[14][23] ),
    .A3(\dpath.RF.R[15][23] ),
    .S0(net569),
    .S1(net550),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_1 _10091_ (.A0(\dpath.RF.R[8][23] ),
    .A1(\dpath.RF.R[9][23] ),
    .A2(\dpath.RF.R[10][23] ),
    .A3(\dpath.RF.R[11][23] ),
    .S0(net569),
    .S1(net550),
    .X(_04286_));
 sky130_fd_sc_hd__or2_1 _10092_ (.A(net534),
    .B(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__o211a_1 _10093_ (.A1(net513),
    .A2(_04285_),
    .B1(_04287_),
    .C1(net528),
    .X(_04288_));
 sky130_fd_sc_hd__nor2_1 _10094_ (.A(net519),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__mux4_1 _10095_ (.A0(\dpath.RF.R[16][23] ),
    .A1(\dpath.RF.R[17][23] ),
    .A2(\dpath.RF.R[18][23] ),
    .A3(\dpath.RF.R[19][23] ),
    .S0(net573),
    .S1(net554),
    .X(_04290_));
 sky130_fd_sc_hd__nor2_1 _10096_ (.A(net536),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__mux4_1 _10097_ (.A0(\dpath.RF.R[20][23] ),
    .A1(\dpath.RF.R[21][23] ),
    .A2(\dpath.RF.R[22][23] ),
    .A3(\dpath.RF.R[23][23] ),
    .S0(net571),
    .S1(net552),
    .X(_04292_));
 sky130_fd_sc_hd__nor2_1 _10098_ (.A(net515),
    .B(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__mux4_1 _10099_ (.A0(\dpath.RF.R[28][23] ),
    .A1(\dpath.RF.R[29][23] ),
    .A2(\dpath.RF.R[30][23] ),
    .A3(\dpath.RF.R[31][23] ),
    .S0(net573),
    .S1(net554),
    .X(_04294_));
 sky130_fd_sc_hd__nor2_1 _10100_ (.A(net515),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__mux4_1 _10101_ (.A0(\dpath.RF.R[24][23] ),
    .A1(\dpath.RF.R[25][23] ),
    .A2(\dpath.RF.R[26][23] ),
    .A3(\dpath.RF.R[27][23] ),
    .S0(net573),
    .S1(net554),
    .X(_04296_));
 sky130_fd_sc_hd__o21ai_1 _10102_ (.A1(net536),
    .A2(_04296_),
    .B1(net526),
    .Y(_04297_));
 sky130_fd_sc_hd__o32a_1 _10103_ (.A1(net526),
    .A2(_04291_),
    .A3(_04293_),
    .B1(_04295_),
    .B2(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__a221o_1 _10104_ (.A1(_04284_),
    .A2(_04289_),
    .B1(_04298_),
    .B2(net519),
    .C1(net483),
    .X(_04299_));
 sky130_fd_sc_hd__nor2_1 _10105_ (.A(net371),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__mux2_2 _10106_ (.A0(net3636),
    .A1(net16),
    .S(net479),
    .X(_04301_));
 sky130_fd_sc_hd__a221o_2 _10107_ (.A1(net671),
    .A2(net369),
    .B1(net367),
    .B2(_04301_),
    .C1(_04300_),
    .X(_04302_));
 sky130_fd_sc_hd__nand4_2 _10108_ (.A(net648),
    .B(net644),
    .C(net724),
    .D(\dpath.alu.adder.in1[22] ),
    .Y(_04303_));
 sky130_fd_sc_hd__a22o_1 _10109_ (.A1(net645),
    .A2(net724),
    .B1(\dpath.alu.adder.in1[22] ),
    .B2(net648),
    .X(_04304_));
 sky130_fd_sc_hd__nand4_2 _10110_ (.A(net639),
    .B(\dpath.alu.adder.in1[20] ),
    .C(_04303_),
    .D(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__a22o_1 _10111_ (.A1(net639),
    .A2(\dpath.alu.adder.in1[20] ),
    .B1(_04303_),
    .B2(_04304_),
    .X(_04306_));
 sky130_fd_sc_hd__o211a_1 _10112_ (.A1(_04196_),
    .A2(_04198_),
    .B1(_04305_),
    .C1(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__a211oi_2 _10113_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_04196_),
    .C1(_04198_),
    .Y(_04308_));
 sky130_fd_sc_hd__nor2_1 _10114_ (.A(_04307_),
    .B(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__and4_1 _10115_ (.A(net635),
    .B(net631),
    .C(\dpath.alu.adder.in1[18] ),
    .D(net727),
    .X(_04310_));
 sky130_fd_sc_hd__a22o_1 _10116_ (.A1(net631),
    .A2(\dpath.alu.adder.in1[18] ),
    .B1(net727),
    .B2(net635),
    .X(_04311_));
 sky130_fd_sc_hd__nand2b_1 _10117_ (.A_N(_04310_),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand2_1 _10118_ (.A(net626),
    .B(net730),
    .Y(_04313_));
 sky130_fd_sc_hd__xnor2_2 _10119_ (.A(_04312_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__xnor2_1 _10120_ (.A(_04309_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__o21ai_2 _10121_ (.A1(_04200_),
    .A2(_04208_),
    .B1(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__or3_1 _10122_ (.A(_04200_),
    .B(_04208_),
    .C(_04315_),
    .X(_04317_));
 sky130_fd_sc_hd__nand4_2 _10123_ (.A(net652),
    .B(\dpath.alu.adder.in1[23] ),
    .C(_04316_),
    .D(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__a22o_1 _10124_ (.A1(net652),
    .A2(net721),
    .B1(_04316_),
    .B2(_04317_),
    .X(_04319_));
 sky130_fd_sc_hd__and2_1 _10125_ (.A(_04318_),
    .B(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__and3_1 _10126_ (.A(net755),
    .B(net752),
    .C(net601),
    .X(_04321_));
 sky130_fd_sc_hd__a22o_1 _10127_ (.A1(net752),
    .A2(net601),
    .B1(net598),
    .B2(net755),
    .X(_04322_));
 sky130_fd_sc_hd__a21bo_1 _10128_ (.A1(net598),
    .A2(_04321_),
    .B1_N(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__nand2_1 _10129_ (.A(net758),
    .B(net596),
    .Y(_04324_));
 sky130_fd_sc_hd__xor2_2 _10130_ (.A(_04323_),
    .B(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__and4_1 _10131_ (.A(net610),
    .B(net607),
    .C(net746),
    .D(net742),
    .X(_04326_));
 sky130_fd_sc_hd__nand4_1 _10132_ (.A(net610),
    .B(net607),
    .C(net746),
    .D(net742),
    .Y(_04327_));
 sky130_fd_sc_hd__a22o_1 _10133_ (.A1(net607),
    .A2(net746),
    .B1(net742),
    .B2(net610),
    .X(_04328_));
 sky130_fd_sc_hd__and4_1 _10134_ (.A(net750),
    .B(net604),
    .C(_04327_),
    .D(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__nand4_1 _10135_ (.A(net750),
    .B(net604),
    .C(_04327_),
    .D(_04328_),
    .Y(_04330_));
 sky130_fd_sc_hd__a22o_1 _10136_ (.A1(net750),
    .A2(net604),
    .B1(_04327_),
    .B2(_04328_),
    .X(_04331_));
 sky130_fd_sc_hd__o211a_1 _10137_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04330_),
    .C1(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__a211o_1 _10138_ (.A1(_04330_),
    .A2(_04331_),
    .B1(_04218_),
    .C1(_04219_),
    .X(_04333_));
 sky130_fd_sc_hd__nand2b_1 _10139_ (.A_N(_04332_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__xnor2_2 _10140_ (.A(_04325_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__nand2_1 _10141_ (.A(_04229_),
    .B(_04231_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand4_2 _10142_ (.A(net623),
    .B(net619),
    .C(\dpath.alu.adder.in1[15] ),
    .D(net733),
    .Y(_04337_));
 sky130_fd_sc_hd__a22o_1 _10143_ (.A1(net619),
    .A2(\dpath.alu.adder.in1[15] ),
    .B1(\dpath.alu.adder.in1[16] ),
    .B2(net622),
    .X(_04338_));
 sky130_fd_sc_hd__nand4_2 _10144_ (.A(net614),
    .B(net737),
    .C(_04337_),
    .D(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__a22o_1 _10145_ (.A1(net615),
    .A2(net737),
    .B1(_04337_),
    .B2(_04338_),
    .X(_04340_));
 sky130_fd_sc_hd__o211ai_2 _10146_ (.A1(_04203_),
    .A2(_04206_),
    .B1(_04339_),
    .C1(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__a211o_1 _10147_ (.A1(_04339_),
    .A2(_04340_),
    .B1(_04203_),
    .C1(_04206_),
    .X(_04342_));
 sky130_fd_sc_hd__nand3_1 _10148_ (.A(_04336_),
    .B(_04341_),
    .C(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__a21o_1 _10149_ (.A1(_04341_),
    .A2(_04342_),
    .B1(_04336_),
    .X(_04344_));
 sky130_fd_sc_hd__a21bo_1 _10150_ (.A1(_04226_),
    .A2(_04233_),
    .B1_N(_04232_),
    .X(_04345_));
 sky130_fd_sc_hd__and3_1 _10151_ (.A(_04343_),
    .B(_04344_),
    .C(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__nand3_1 _10152_ (.A(_04343_),
    .B(_04344_),
    .C(_04345_),
    .Y(_04347_));
 sky130_fd_sc_hd__a21o_1 _10153_ (.A1(_04343_),
    .A2(_04344_),
    .B1(_04345_),
    .X(_04348_));
 sky130_fd_sc_hd__and3_2 _10154_ (.A(_04335_),
    .B(_04347_),
    .C(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__a21oi_1 _10155_ (.A1(_04347_),
    .A2(_04348_),
    .B1(_04335_),
    .Y(_04350_));
 sky130_fd_sc_hd__or3_2 _10156_ (.A(_04210_),
    .B(_04349_),
    .C(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__o21ai_2 _10157_ (.A1(_04349_),
    .A2(_04350_),
    .B1(_04210_),
    .Y(_04352_));
 sky130_fd_sc_hd__o211ai_4 _10158_ (.A1(_04237_),
    .A2(_04240_),
    .B1(_04351_),
    .C1(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__a211o_1 _10159_ (.A1(_04351_),
    .A2(_04352_),
    .B1(_04237_),
    .C1(_04240_),
    .X(_04354_));
 sky130_fd_sc_hd__and3_1 _10160_ (.A(_04320_),
    .B(_04353_),
    .C(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__a21oi_1 _10161_ (.A1(_04353_),
    .A2(_04354_),
    .B1(_04320_),
    .Y(_04356_));
 sky130_fd_sc_hd__o21a_1 _10162_ (.A1(_04355_),
    .A2(_04356_),
    .B1(_04246_),
    .X(_04357_));
 sky130_fd_sc_hd__nor3_1 _10163_ (.A(_04246_),
    .B(_04355_),
    .C(_04356_),
    .Y(_04358_));
 sky130_fd_sc_hd__or3_2 _10164_ (.A(_04246_),
    .B(_04355_),
    .C(_04356_),
    .X(_04359_));
 sky130_fd_sc_hd__a22oi_1 _10165_ (.A1(net773),
    .A2(net586),
    .B1(net584),
    .B2(net778),
    .Y(_04360_));
 sky130_fd_sc_hd__and4_1 _10166_ (.A(net778),
    .B(net773),
    .C(net586),
    .D(net584),
    .X(_04361_));
 sky130_fd_sc_hd__o2bb2a_1 _10167_ (.A1_N(net782),
    .A2_N(net582),
    .B1(_04360_),
    .B2(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__and4bb_1 _10168_ (.A_N(_04360_),
    .B_N(_04361_),
    .C(net782),
    .D(net582),
    .X(_04363_));
 sky130_fd_sc_hd__or2_1 _10169_ (.A(_04362_),
    .B(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__or2_2 _10170_ (.A(_04156_),
    .B(_04158_),
    .X(_04365_));
 sky130_fd_sc_hd__and2b_1 _10171_ (.A_N(_04364_),
    .B(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__xnor2_2 _10172_ (.A(_04364_),
    .B(_04365_),
    .Y(_04367_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(\dpath.alu.adder.in1[1] ),
    .B(net580),
    .Y(_04368_));
 sky130_fd_sc_hd__inv_2 _10174_ (.A(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__xnor2_1 _10175_ (.A(_04367_),
    .B(_04368_),
    .Y(_04370_));
 sky130_fd_sc_hd__a31o_1 _10176_ (.A1(net785),
    .A2(net582),
    .A3(_04162_),
    .B1(_04161_),
    .X(_04371_));
 sky130_fd_sc_hd__xor2_1 _10177_ (.A(_04370_),
    .B(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _10178_ (.A(net789),
    .B(\dpath.alu.adder.in0[23] ),
    .Y(_04373_));
 sky130_fd_sc_hd__and3_1 _10179_ (.A(\dpath.alu.adder.in1[0] ),
    .B(\dpath.alu.adder.in0[23] ),
    .C(_04372_),
    .X(_04374_));
 sky130_fd_sc_hd__xor2_1 _10180_ (.A(_04372_),
    .B(_04373_),
    .X(_04375_));
 sky130_fd_sc_hd__a31o_1 _10181_ (.A1(_04214_),
    .A2(_04215_),
    .A3(_04223_),
    .B1(_04222_),
    .X(_04376_));
 sky130_fd_sc_hd__nand2_1 _10182_ (.A(_04175_),
    .B(_04177_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand4_1 _10183_ (.A(net766),
    .B(net760),
    .C(net593),
    .D(net590),
    .Y(_04378_));
 sky130_fd_sc_hd__a22o_1 _10184_ (.A1(net760),
    .A2(net593),
    .B1(net590),
    .B2(net766),
    .X(_04379_));
 sky130_fd_sc_hd__and4_1 _10185_ (.A(net769),
    .B(net587),
    .C(_04378_),
    .D(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__a22oi_2 _10186_ (.A1(net769),
    .A2(net588),
    .B1(_04378_),
    .B2(_04379_),
    .Y(_04381_));
 sky130_fd_sc_hd__a211o_2 _10187_ (.A1(_04213_),
    .A2(_04215_),
    .B1(_04380_),
    .C1(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__o211ai_2 _10188_ (.A1(_04380_),
    .A2(_04381_),
    .B1(_04213_),
    .C1(_04215_),
    .Y(_04383_));
 sky130_fd_sc_hd__nand3_2 _10189_ (.A(_04377_),
    .B(_04382_),
    .C(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a21o_1 _10190_ (.A1(_04382_),
    .A2(_04383_),
    .B1(_04377_),
    .X(_04385_));
 sky130_fd_sc_hd__and3_2 _10191_ (.A(_04376_),
    .B(_04384_),
    .C(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__a21oi_2 _10192_ (.A1(_04384_),
    .A2(_04385_),
    .B1(_04376_),
    .Y(_04387_));
 sky130_fd_sc_hd__a211oi_4 _10193_ (.A1(_04178_),
    .A2(_04180_),
    .B1(_04386_),
    .C1(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__o211a_1 _10194_ (.A1(_04386_),
    .A2(_04387_),
    .B1(_04178_),
    .C1(_04180_),
    .X(_04389_));
 sky130_fd_sc_hd__a211oi_4 _10195_ (.A1(_04183_),
    .A2(_04185_),
    .B1(_04388_),
    .C1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__inv_2 _10196_ (.A(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__o211a_1 _10197_ (.A1(_04388_),
    .A2(_04389_),
    .B1(_04183_),
    .C1(_04185_),
    .X(_04392_));
 sky130_fd_sc_hd__nor3_2 _10198_ (.A(_04375_),
    .B(_04390_),
    .C(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__inv_2 _10199_ (.A(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__o21a_1 _10200_ (.A1(_04390_),
    .A2(_04392_),
    .B1(_04375_),
    .X(_04395_));
 sky130_fd_sc_hd__a211o_1 _10201_ (.A1(_04242_),
    .A2(_04244_),
    .B1(_04393_),
    .C1(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__o211ai_2 _10202_ (.A1(_04393_),
    .A2(_04395_),
    .B1(_04242_),
    .C1(_04244_),
    .Y(_04397_));
 sky130_fd_sc_hd__o211a_1 _10203_ (.A1(_04187_),
    .A2(_04189_),
    .B1(_04396_),
    .C1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__inv_2 _10204_ (.A(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__a211oi_2 _10205_ (.A1(_04396_),
    .A2(_04397_),
    .B1(_04187_),
    .C1(_04189_),
    .Y(_04400_));
 sky130_fd_sc_hd__or4_4 _10206_ (.A(_04357_),
    .B(_04358_),
    .C(_04398_),
    .D(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__o22ai_2 _10207_ (.A1(_04357_),
    .A2(_04358_),
    .B1(_04398_),
    .B2(_04400_),
    .Y(_04402_));
 sky130_fd_sc_hd__o211a_1 _10208_ (.A1(_04249_),
    .A2(_04251_),
    .B1(_04401_),
    .C1(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__a211oi_2 _10209_ (.A1(_04401_),
    .A2(_04402_),
    .B1(_04249_),
    .C1(_04251_),
    .Y(_04404_));
 sky130_fd_sc_hd__a211oi_2 _10210_ (.A1(_04191_),
    .A2(_04193_),
    .B1(_04403_),
    .C1(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__o211a_1 _10211_ (.A1(_04403_),
    .A2(_04404_),
    .B1(_04191_),
    .C1(_04193_),
    .X(_04406_));
 sky130_fd_sc_hd__a211oi_2 _10212_ (.A1(_04254_),
    .A2(_04256_),
    .B1(_04405_),
    .C1(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__o211a_1 _10213_ (.A1(_04405_),
    .A2(_04406_),
    .B1(_04254_),
    .C1(_04256_),
    .X(_04408_));
 sky130_fd_sc_hd__a211oi_2 _10214_ (.A1(_04166_),
    .A2(_04169_),
    .B1(_04407_),
    .C1(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__o211a_1 _10215_ (.A1(_04407_),
    .A2(_04408_),
    .B1(_04166_),
    .C1(_04169_),
    .X(_04410_));
 sky130_fd_sc_hd__o211a_1 _10216_ (.A1(_04409_),
    .A2(_04410_),
    .B1(_04258_),
    .C1(_04261_),
    .X(_04411_));
 sky130_fd_sc_hd__a211oi_2 _10217_ (.A1(_04258_),
    .A2(_04261_),
    .B1(_04409_),
    .C1(_04410_),
    .Y(_04412_));
 sky130_fd_sc_hd__nor2_1 _10218_ (.A(_04411_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21ai_1 _10219_ (.A1(_04263_),
    .A2(_04270_),
    .B1(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__or3_1 _10220_ (.A(_04263_),
    .B(_04270_),
    .C(_04413_),
    .X(_04415_));
 sky130_fd_sc_hd__a21o_1 _10221_ (.A1(_04414_),
    .A2(_04415_),
    .B1(net486),
    .X(_04416_));
 sky130_fd_sc_hd__o21a_1 _10222_ (.A1(net3626),
    .A2(_02071_),
    .B1(net469),
    .X(_04417_));
 sky130_fd_sc_hd__a21oi_1 _10223_ (.A1(_01921_),
    .A2(_04272_),
    .B1(_01919_),
    .Y(_04418_));
 sky130_fd_sc_hd__a31o_1 _10224_ (.A1(_01919_),
    .A2(_01921_),
    .A3(_04272_),
    .B1(net469),
    .X(_04419_));
 sky130_fd_sc_hd__nor2_1 _10225_ (.A(_04418_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__a21o_4 _10226_ (.A1(_04416_),
    .A2(_04417_),
    .B1(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__a21oi_4 _10227_ (.A1(net391),
    .A2(_04421_),
    .B1(_04302_),
    .Y(_04422_));
 sky130_fd_sc_hd__xnor2_1 _10228_ (.A(net577),
    .B(net3468),
    .Y(_04423_));
 sky130_fd_sc_hd__a21o_1 _10229_ (.A1(net577),
    .A2(net3466),
    .B1(_04127_),
    .X(_04424_));
 sky130_fd_sc_hd__xor2_1 _10230_ (.A(_04423_),
    .B(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__and2_1 _10231_ (.A(net3546),
    .B(_04278_),
    .X(_04426_));
 sky130_fd_sc_hd__nor2_1 _10232_ (.A(net3546),
    .B(_04278_),
    .Y(_04427_));
 sky130_fd_sc_hd__or3_1 _10233_ (.A(_01958_),
    .B(_04426_),
    .C(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__a21oi_1 _10234_ (.A1(\dpath.btarg_DX.q[23] ),
    .A2(net404),
    .B1(net452),
    .Y(_04429_));
 sky130_fd_sc_hd__o211a_1 _10235_ (.A1(net366),
    .A2(_04425_),
    .B1(_04428_),
    .C1(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__o21ai_1 _10236_ (.A1(net374),
    .A2(_04422_),
    .B1(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__o211a_1 _10237_ (.A1(net3546),
    .A2(net445),
    .B1(_04431_),
    .C1(net851),
    .X(_00659_));
 sky130_fd_sc_hd__mux4_1 _10238_ (.A0(\dpath.RF.R[0][24] ),
    .A1(\dpath.RF.R[1][24] ),
    .A2(\dpath.RF.R[2][24] ),
    .A3(\dpath.RF.R[3][24] ),
    .S0(net569),
    .S1(net550),
    .X(_04432_));
 sky130_fd_sc_hd__mux4_1 _10239_ (.A0(\dpath.RF.R[4][24] ),
    .A1(\dpath.RF.R[5][24] ),
    .A2(\dpath.RF.R[6][24] ),
    .A3(\dpath.RF.R[7][24] ),
    .S0(net569),
    .S1(net550),
    .X(_04433_));
 sky130_fd_sc_hd__o21a_1 _10240_ (.A1(net514),
    .A2(_04433_),
    .B1(net507),
    .X(_04434_));
 sky130_fd_sc_hd__o21ai_1 _10241_ (.A1(net534),
    .A2(_04432_),
    .B1(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__mux4_1 _10242_ (.A0(\dpath.RF.R[12][24] ),
    .A1(\dpath.RF.R[13][24] ),
    .A2(\dpath.RF.R[14][24] ),
    .A3(\dpath.RF.R[15][24] ),
    .S0(net569),
    .S1(net550),
    .X(_04436_));
 sky130_fd_sc_hd__mux4_1 _10243_ (.A0(\dpath.RF.R[8][24] ),
    .A1(\dpath.RF.R[9][24] ),
    .A2(\dpath.RF.R[10][24] ),
    .A3(\dpath.RF.R[11][24] ),
    .S0(net569),
    .S1(net550),
    .X(_04437_));
 sky130_fd_sc_hd__or2_1 _10244_ (.A(net534),
    .B(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__o211a_1 _10245_ (.A1(net513),
    .A2(_04436_),
    .B1(_04438_),
    .C1(net528),
    .X(_04439_));
 sky130_fd_sc_hd__nor2_1 _10246_ (.A(net519),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__mux4_1 _10247_ (.A0(\dpath.RF.R[16][24] ),
    .A1(\dpath.RF.R[17][24] ),
    .A2(\dpath.RF.R[18][24] ),
    .A3(\dpath.RF.R[19][24] ),
    .S0(net570),
    .S1(net551),
    .X(_04441_));
 sky130_fd_sc_hd__nor2_1 _10248_ (.A(_00007_),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__mux4_1 _10249_ (.A0(\dpath.RF.R[20][24] ),
    .A1(\dpath.RF.R[21][24] ),
    .A2(\dpath.RF.R[22][24] ),
    .A3(\dpath.RF.R[23][24] ),
    .S0(net569),
    .S1(net550),
    .X(_04443_));
 sky130_fd_sc_hd__nor2_1 _10250_ (.A(net513),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__mux4_1 _10251_ (.A0(\dpath.RF.R[28][24] ),
    .A1(\dpath.RF.R[29][24] ),
    .A2(\dpath.RF.R[30][24] ),
    .A3(\dpath.RF.R[31][24] ),
    .S0(net570),
    .S1(net551),
    .X(_04445_));
 sky130_fd_sc_hd__nor2_1 _10252_ (.A(_01771_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__mux4_1 _10253_ (.A0(\dpath.RF.R[24][24] ),
    .A1(\dpath.RF.R[25][24] ),
    .A2(\dpath.RF.R[26][24] ),
    .A3(\dpath.RF.R[27][24] ),
    .S0(net569),
    .S1(net550),
    .X(_04447_));
 sky130_fd_sc_hd__o21ai_1 _10254_ (.A1(_00007_),
    .A2(_04447_),
    .B1(net528),
    .Y(_04448_));
 sky130_fd_sc_hd__o32a_1 _10255_ (.A1(net528),
    .A2(_04442_),
    .A3(_04444_),
    .B1(_04446_),
    .B2(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__a221o_1 _10256_ (.A1(_04435_),
    .A2(_04440_),
    .B1(_04449_),
    .B2(net519),
    .C1(net483),
    .X(_04450_));
 sky130_fd_sc_hd__nor2_1 _10257_ (.A(net371),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__mux2_2 _10258_ (.A0(net3632),
    .A1(net17),
    .S(net479),
    .X(_04452_));
 sky130_fd_sc_hd__a221o_2 _10259_ (.A1(net670),
    .A2(net369),
    .B1(net367),
    .B2(_04452_),
    .C1(_04451_),
    .X(_04453_));
 sky130_fd_sc_hd__a31o_1 _10260_ (.A1(_01918_),
    .A2(_01921_),
    .A3(_04272_),
    .B1(_01917_),
    .X(_04454_));
 sky130_fd_sc_hd__nand2_1 _10261_ (.A(_01900_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__or2_1 _10262_ (.A(_01900_),
    .B(_04454_),
    .X(_04456_));
 sky130_fd_sc_hd__or4_1 _10263_ (.A(_04263_),
    .B(_04264_),
    .C(_04411_),
    .D(_04412_),
    .X(_04457_));
 sky130_fd_sc_hd__a211o_1 _10264_ (.A1(_03959_),
    .A2(_03960_),
    .B1(_04267_),
    .C1(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__nor2_1 _10265_ (.A(_04266_),
    .B(_04457_),
    .Y(_04459_));
 sky130_fd_sc_hd__and2b_1 _10266_ (.A_N(_04411_),
    .B(_04263_),
    .X(_04460_));
 sky130_fd_sc_hd__nor3_1 _10267_ (.A(_04412_),
    .B(_04459_),
    .C(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__and2_1 _10268_ (.A(_04458_),
    .B(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__a21oi_1 _10269_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04374_),
    .Y(_04463_));
 sky130_fd_sc_hd__a22o_1 _10270_ (.A1(net648),
    .A2(\dpath.alu.adder.in1[23] ),
    .B1(net720),
    .B2(net652),
    .X(_04464_));
 sky130_fd_sc_hd__and3_1 _10271_ (.A(net652),
    .B(net648),
    .C(net720),
    .X(_04465_));
 sky130_fd_sc_hd__and2_1 _10272_ (.A(net721),
    .B(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(\dpath.alu.adder.in1[23] ),
    .B(_04465_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _10274_ (.A(_04464_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__and4_1 _10275_ (.A(net644),
    .B(net640),
    .C(net723),
    .D(net722),
    .X(_04469_));
 sky130_fd_sc_hd__a22o_1 _10276_ (.A1(net640),
    .A2(net723),
    .B1(\dpath.alu.adder.in1[22] ),
    .B2(net644),
    .X(_04470_));
 sky130_fd_sc_hd__nand2b_1 _10277_ (.A_N(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(net634),
    .B(\dpath.alu.adder.in1[20] ),
    .Y(_04472_));
 sky130_fd_sc_hd__xnor2_2 _10279_ (.A(_04471_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__nand2_1 _10280_ (.A(_04303_),
    .B(_04305_),
    .Y(_04474_));
 sky130_fd_sc_hd__and2b_1 _10281_ (.A_N(_04473_),
    .B(_04474_),
    .X(_04475_));
 sky130_fd_sc_hd__xor2_2 _10282_ (.A(_04473_),
    .B(_04474_),
    .X(_04476_));
 sky130_fd_sc_hd__nand4_1 _10283_ (.A(net630),
    .B(net626),
    .C(net729),
    .D(net726),
    .Y(_04477_));
 sky130_fd_sc_hd__a22o_1 _10284_ (.A1(net626),
    .A2(net729),
    .B1(net726),
    .B2(net630),
    .X(_04478_));
 sky130_fd_sc_hd__nand2_1 _10285_ (.A(_04477_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__and2_1 _10286_ (.A(net622),
    .B(net730),
    .X(_04480_));
 sky130_fd_sc_hd__xor2_2 _10287_ (.A(_04479_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__nor2_1 _10288_ (.A(_04476_),
    .B(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__xor2_2 _10289_ (.A(_04476_),
    .B(_04481_),
    .X(_04483_));
 sky130_fd_sc_hd__o21bai_2 _10290_ (.A1(_04308_),
    .A2(_04314_),
    .B1_N(_04307_),
    .Y(_04484_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_04483_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__xor2_2 _10292_ (.A(_04483_),
    .B(_04484_),
    .X(_04486_));
 sky130_fd_sc_hd__and3_1 _10293_ (.A(_04464_),
    .B(_04467_),
    .C(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__xor2_2 _10294_ (.A(_04468_),
    .B(_04486_),
    .X(_04488_));
 sky130_fd_sc_hd__nor2_2 _10295_ (.A(_04318_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__xor2_1 _10296_ (.A(_04318_),
    .B(_04488_),
    .X(_04490_));
 sky130_fd_sc_hd__and3_1 _10297_ (.A(net756),
    .B(net753),
    .C(net598),
    .X(_04491_));
 sky130_fd_sc_hd__a22o_1 _10298_ (.A1(net753),
    .A2(net598),
    .B1(net596),
    .B2(net756),
    .X(_04492_));
 sky130_fd_sc_hd__a21bo_1 _10299_ (.A1(net596),
    .A2(_04491_),
    .B1_N(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__nand2_1 _10300_ (.A(net759),
    .B(net592),
    .Y(_04494_));
 sky130_fd_sc_hd__xor2_2 _10301_ (.A(_04493_),
    .B(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__a22o_1 _10302_ (.A1(net604),
    .A2(net746),
    .B1(net742),
    .B2(net607),
    .X(_04496_));
 sky130_fd_sc_hd__and4_1 _10303_ (.A(net607),
    .B(net604),
    .C(net743),
    .D(net739),
    .X(_04497_));
 sky130_fd_sc_hd__nand4_1 _10304_ (.A(net607),
    .B(net604),
    .C(net746),
    .D(net742),
    .Y(_04498_));
 sky130_fd_sc_hd__and4_1 _10305_ (.A(net747),
    .B(net601),
    .C(_04496_),
    .D(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__nand4_1 _10306_ (.A(net750),
    .B(net601),
    .C(_04496_),
    .D(_04498_),
    .Y(_04500_));
 sky130_fd_sc_hd__a22o_1 _10307_ (.A1(net750),
    .A2(net601),
    .B1(_04496_),
    .B2(_04498_),
    .X(_04501_));
 sky130_fd_sc_hd__o211a_1 _10308_ (.A1(_04326_),
    .A2(_04329_),
    .B1(_04500_),
    .C1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__a211o_1 _10309_ (.A1(_04500_),
    .A2(_04501_),
    .B1(_04326_),
    .C1(_04329_),
    .X(_04503_));
 sky130_fd_sc_hd__nand2b_1 _10310_ (.A_N(_04502_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__xnor2_2 _10311_ (.A(_04495_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__nand2_1 _10312_ (.A(_04337_),
    .B(_04339_),
    .Y(_04506_));
 sky130_fd_sc_hd__a31o_1 _10313_ (.A1(net627),
    .A2(net730),
    .A3(_04311_),
    .B1(_04310_),
    .X(_04507_));
 sky130_fd_sc_hd__nand4_2 _10314_ (.A(net618),
    .B(net614),
    .C(\dpath.alu.adder.in1[15] ),
    .D(\dpath.alu.adder.in1[16] ),
    .Y(_04508_));
 sky130_fd_sc_hd__a22o_1 _10315_ (.A1(net614),
    .A2(\dpath.alu.adder.in1[15] ),
    .B1(\dpath.alu.adder.in1[16] ),
    .B2(net618),
    .X(_04509_));
 sky130_fd_sc_hd__nand4_2 _10316_ (.A(net610),
    .B(net737),
    .C(_04508_),
    .D(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__a22o_1 _10317_ (.A1(net610),
    .A2(net737),
    .B1(_04508_),
    .B2(_04509_),
    .X(_04511_));
 sky130_fd_sc_hd__nand3_1 _10318_ (.A(_04507_),
    .B(_04510_),
    .C(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__a21o_1 _10319_ (.A1(_04510_),
    .A2(_04511_),
    .B1(_04507_),
    .X(_04513_));
 sky130_fd_sc_hd__nand3_1 _10320_ (.A(_04506_),
    .B(_04512_),
    .C(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__a21o_1 _10321_ (.A1(_04512_),
    .A2(_04513_),
    .B1(_04506_),
    .X(_04515_));
 sky130_fd_sc_hd__a21bo_1 _10322_ (.A1(_04336_),
    .A2(_04342_),
    .B1_N(_04341_),
    .X(_04516_));
 sky130_fd_sc_hd__and3_1 _10323_ (.A(_04514_),
    .B(_04515_),
    .C(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__nand3_1 _10324_ (.A(_04514_),
    .B(_04515_),
    .C(_04516_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21o_1 _10325_ (.A1(_04514_),
    .A2(_04515_),
    .B1(_04516_),
    .X(_04519_));
 sky130_fd_sc_hd__and3_2 _10326_ (.A(_04505_),
    .B(_04518_),
    .C(_04519_),
    .X(_04520_));
 sky130_fd_sc_hd__a21oi_1 _10327_ (.A1(_04518_),
    .A2(_04519_),
    .B1(_04505_),
    .Y(_04521_));
 sky130_fd_sc_hd__or3_4 _10328_ (.A(_04316_),
    .B(_04520_),
    .C(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__o21ai_2 _10329_ (.A1(_04520_),
    .A2(_04521_),
    .B1(_04316_),
    .Y(_04523_));
 sky130_fd_sc_hd__o211ai_4 _10330_ (.A1(_04346_),
    .A2(_04349_),
    .B1(_04522_),
    .C1(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__a211o_1 _10331_ (.A1(_04522_),
    .A2(_04523_),
    .B1(_04346_),
    .C1(_04349_),
    .X(_04525_));
 sky130_fd_sc_hd__and3_2 _10332_ (.A(_04490_),
    .B(_04524_),
    .C(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__nand3_1 _10333_ (.A(_04490_),
    .B(_04524_),
    .C(_04525_),
    .Y(_04527_));
 sky130_fd_sc_hd__a21o_1 _10334_ (.A1(_04524_),
    .A2(_04525_),
    .B1(_04490_),
    .X(_04528_));
 sky130_fd_sc_hd__a21oi_2 _10335_ (.A1(_04527_),
    .A2(_04528_),
    .B1(_04355_),
    .Y(_04529_));
 sky130_fd_sc_hd__and3_1 _10336_ (.A(_04355_),
    .B(_04527_),
    .C(_04528_),
    .X(_04530_));
 sky130_fd_sc_hd__inv_2 _10337_ (.A(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__and4_1 _10338_ (.A(net777),
    .B(net773),
    .C(net584),
    .D(net582),
    .X(_04532_));
 sky130_fd_sc_hd__a22o_1 _10339_ (.A1(net773),
    .A2(net584),
    .B1(net582),
    .B2(net777),
    .X(_04533_));
 sky130_fd_sc_hd__nand2b_1 _10340_ (.A_N(_04532_),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _10341_ (.A(net782),
    .B(net580),
    .Y(_04535_));
 sky130_fd_sc_hd__xnor2_2 _10342_ (.A(_04534_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__or2_1 _10343_ (.A(_04361_),
    .B(_04363_),
    .X(_04537_));
 sky130_fd_sc_hd__and2b_1 _10344_ (.A_N(_04536_),
    .B(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__xnor2_2 _10345_ (.A(_04536_),
    .B(_04537_),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _10346_ (.A(net784),
    .B(net579),
    .Y(_04540_));
 sky130_fd_sc_hd__xor2_2 _10347_ (.A(_04539_),
    .B(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__a21oi_2 _10348_ (.A1(_04367_),
    .A2(_04369_),
    .B1(_04366_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_1 _10349_ (.A(_04541_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__xor2_2 _10350_ (.A(_04541_),
    .B(_04542_),
    .X(_04544_));
 sky130_fd_sc_hd__nand2_1 _10351_ (.A(net789),
    .B(\dpath.alu.adder.in0[24] ),
    .Y(_04545_));
 sky130_fd_sc_hd__xor2_2 _10352_ (.A(_04544_),
    .B(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__a21o_1 _10353_ (.A1(_04325_),
    .A2(_04333_),
    .B1(_04332_),
    .X(_04547_));
 sky130_fd_sc_hd__a41o_1 _10354_ (.A1(net764),
    .A2(net763),
    .A3(net593),
    .A4(net590),
    .B1(_04380_),
    .X(_04548_));
 sky130_fd_sc_hd__a32o_1 _10355_ (.A1(net758),
    .A2(net596),
    .A3(_04322_),
    .B1(_04321_),
    .B2(net599),
    .X(_04549_));
 sky130_fd_sc_hd__nand4_2 _10356_ (.A(net764),
    .B(net760),
    .C(net590),
    .D(net588),
    .Y(_04550_));
 sky130_fd_sc_hd__a22o_1 _10357_ (.A1(net760),
    .A2(net590),
    .B1(net588),
    .B2(\dpath.alu.adder.in1[6] ),
    .X(_04551_));
 sky130_fd_sc_hd__nand4_2 _10358_ (.A(net771),
    .B(net585),
    .C(_04550_),
    .D(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a22o_1 _10359_ (.A1(net768),
    .A2(net586),
    .B1(_04550_),
    .B2(_04551_),
    .X(_04553_));
 sky130_fd_sc_hd__nand3_2 _10360_ (.A(_04549_),
    .B(_04552_),
    .C(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__a21o_1 _10361_ (.A1(_04552_),
    .A2(_04553_),
    .B1(_04549_),
    .X(_04555_));
 sky130_fd_sc_hd__nand3_2 _10362_ (.A(_04548_),
    .B(_04554_),
    .C(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__a21o_1 _10363_ (.A1(_04554_),
    .A2(_04555_),
    .B1(_04548_),
    .X(_04557_));
 sky130_fd_sc_hd__and3_2 _10364_ (.A(_04547_),
    .B(_04556_),
    .C(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__a21oi_2 _10365_ (.A1(_04556_),
    .A2(_04557_),
    .B1(_04547_),
    .Y(_04559_));
 sky130_fd_sc_hd__a211oi_1 _10366_ (.A1(_04382_),
    .A2(_04384_),
    .B1(_04558_),
    .C1(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__a211o_1 _10367_ (.A1(_04382_),
    .A2(_04384_),
    .B1(_04558_),
    .C1(_04559_),
    .X(_04561_));
 sky130_fd_sc_hd__o211ai_2 _10368_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04382_),
    .C1(_04384_),
    .Y(_04562_));
 sky130_fd_sc_hd__o211a_2 _10369_ (.A1(_04386_),
    .A2(_04388_),
    .B1(_04561_),
    .C1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__inv_2 _10370_ (.A(_04563_),
    .Y(_04564_));
 sky130_fd_sc_hd__a211oi_2 _10371_ (.A1(_04561_),
    .A2(_04562_),
    .B1(_04386_),
    .C1(_04388_),
    .Y(_04565_));
 sky130_fd_sc_hd__nor3_1 _10372_ (.A(_04546_),
    .B(_04563_),
    .C(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__or3_2 _10373_ (.A(_04546_),
    .B(_04563_),
    .C(_04565_),
    .X(_04567_));
 sky130_fd_sc_hd__o21a_1 _10374_ (.A1(_04563_),
    .A2(_04565_),
    .B1(_04546_),
    .X(_04568_));
 sky130_fd_sc_hd__a211oi_2 _10375_ (.A1(_04351_),
    .A2(_04353_),
    .B1(_04566_),
    .C1(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__o211a_1 _10376_ (.A1(_04566_),
    .A2(_04568_),
    .B1(_04351_),
    .C1(_04353_),
    .X(_04570_));
 sky130_fd_sc_hd__a211oi_2 _10377_ (.A1(_04391_),
    .A2(_04394_),
    .B1(_04569_),
    .C1(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__o211a_1 _10378_ (.A1(_04569_),
    .A2(_04570_),
    .B1(_04391_),
    .C1(_04394_),
    .X(_04572_));
 sky130_fd_sc_hd__nor4_2 _10379_ (.A(_04529_),
    .B(_04530_),
    .C(_04571_),
    .D(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__or4_1 _10380_ (.A(_04529_),
    .B(_04530_),
    .C(_04571_),
    .D(_04572_),
    .X(_04574_));
 sky130_fd_sc_hd__o22a_1 _10381_ (.A1(_04529_),
    .A2(_04530_),
    .B1(_04571_),
    .B2(_04572_),
    .X(_04575_));
 sky130_fd_sc_hd__a211oi_4 _10382_ (.A1(_04359_),
    .A2(_04401_),
    .B1(_04573_),
    .C1(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__o211a_1 _10383_ (.A1(_04573_),
    .A2(_04575_),
    .B1(_04359_),
    .C1(_04401_),
    .X(_04577_));
 sky130_fd_sc_hd__a211oi_2 _10384_ (.A1(_04396_),
    .A2(_04399_),
    .B1(_04576_),
    .C1(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__o211a_1 _10385_ (.A1(_04576_),
    .A2(_04577_),
    .B1(_04396_),
    .C1(_04399_),
    .X(_04579_));
 sky130_fd_sc_hd__nor2_1 _10386_ (.A(_04403_),
    .B(_04405_),
    .Y(_04580_));
 sky130_fd_sc_hd__nor3_2 _10387_ (.A(_04578_),
    .B(_04579_),
    .C(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__o21a_1 _10388_ (.A1(_04578_),
    .A2(_04579_),
    .B1(_04580_),
    .X(_04582_));
 sky130_fd_sc_hd__nor3_1 _10389_ (.A(_04463_),
    .B(_04581_),
    .C(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__o21a_1 _10390_ (.A1(_04581_),
    .A2(_04582_),
    .B1(_04463_),
    .X(_04584_));
 sky130_fd_sc_hd__or2_1 _10391_ (.A(_04583_),
    .B(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__nor2_1 _10392_ (.A(_04407_),
    .B(_04409_),
    .Y(_04586_));
 sky130_fd_sc_hd__nor2_1 _10393_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__xor2_1 _10394_ (.A(_04585_),
    .B(_04586_),
    .X(_04588_));
 sky130_fd_sc_hd__nand2b_1 _10395_ (.A_N(_04588_),
    .B(_04462_),
    .Y(_04589_));
 sky130_fd_sc_hd__and2b_1 _10396_ (.A_N(_04462_),
    .B(_04588_),
    .X(_04590_));
 sky130_fd_sc_hd__nor2_1 _10397_ (.A(_02240_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a32o_1 _10398_ (.A1(net467),
    .A2(_04455_),
    .A3(_04456_),
    .B1(net486),
    .B2(net3687),
    .X(_04592_));
 sky130_fd_sc_hd__a21o_2 _10399_ (.A1(_04589_),
    .A2(_04591_),
    .B1(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__a21o_2 _10400_ (.A1(net391),
    .A2(_04593_),
    .B1(_04453_),
    .X(_04594_));
 sky130_fd_sc_hd__or3_1 _10401_ (.A(_04123_),
    .B(_04125_),
    .C(_04423_),
    .X(_04595_));
 sky130_fd_sc_hd__o41a_1 _10402_ (.A1(net3468),
    .A2(net3466),
    .A3(net3455),
    .A4(net3462),
    .B1(net577),
    .X(_04596_));
 sky130_fd_sc_hd__o21ba_1 _10403_ (.A1(_03975_),
    .A2(_04595_),
    .B1_N(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__or2_1 _10404_ (.A(net577),
    .B(net3542),
    .X(_04598_));
 sky130_fd_sc_hd__nand2_1 _10405_ (.A(net577),
    .B(net3542),
    .Y(_04599_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(_04598_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__xnor2_1 _10407_ (.A(_04597_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__nor2_1 _10408_ (.A(net366),
    .B(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(net3394),
    .B(_04426_),
    .Y(_04603_));
 sky130_fd_sc_hd__o211a_1 _10410_ (.A1(net3394),
    .A2(_04426_),
    .B1(_04603_),
    .C1(net362),
    .X(_04604_));
 sky130_fd_sc_hd__a211o_1 _10411_ (.A1(\dpath.btarg_DX.q[24] ),
    .A2(net404),
    .B1(net452),
    .C1(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__a211o_1 _10412_ (.A1(_02027_),
    .A2(_04594_),
    .B1(_04602_),
    .C1(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o211a_1 _10413_ (.A1(net3394),
    .A2(net445),
    .B1(_04606_),
    .C1(net851),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_1 _10414_ (.A0(\dpath.RF.R[0][25] ),
    .A1(\dpath.RF.R[1][25] ),
    .A2(\dpath.RF.R[2][25] ),
    .A3(\dpath.RF.R[3][25] ),
    .S0(net569),
    .S1(net550),
    .X(_04607_));
 sky130_fd_sc_hd__mux4_1 _10415_ (.A0(\dpath.RF.R[4][25] ),
    .A1(\dpath.RF.R[5][25] ),
    .A2(\dpath.RF.R[6][25] ),
    .A3(\dpath.RF.R[7][25] ),
    .S0(net569),
    .S1(net550),
    .X(_04608_));
 sky130_fd_sc_hd__o21a_1 _10416_ (.A1(_01771_),
    .A2(_04608_),
    .B1(net507),
    .X(_04609_));
 sky130_fd_sc_hd__o21ai_1 _10417_ (.A1(_00007_),
    .A2(_04607_),
    .B1(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__mux4_1 _10418_ (.A0(\dpath.RF.R[12][25] ),
    .A1(\dpath.RF.R[13][25] ),
    .A2(\dpath.RF.R[14][25] ),
    .A3(\dpath.RF.R[15][25] ),
    .S0(net573),
    .S1(net554),
    .X(_04611_));
 sky130_fd_sc_hd__mux4_1 _10419_ (.A0(\dpath.RF.R[8][25] ),
    .A1(\dpath.RF.R[9][25] ),
    .A2(\dpath.RF.R[10][25] ),
    .A3(\dpath.RF.R[11][25] ),
    .S0(net573),
    .S1(net554),
    .X(_04612_));
 sky130_fd_sc_hd__or2_1 _10420_ (.A(net536),
    .B(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__o211a_1 _10421_ (.A1(net515),
    .A2(_04611_),
    .B1(_04613_),
    .C1(net526),
    .X(_04614_));
 sky130_fd_sc_hd__nor2_1 _10422_ (.A(net520),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__mux4_1 _10423_ (.A0(\dpath.RF.R[16][25] ),
    .A1(\dpath.RF.R[17][25] ),
    .A2(\dpath.RF.R[18][25] ),
    .A3(\dpath.RF.R[19][25] ),
    .S0(net573),
    .S1(net554),
    .X(_04616_));
 sky130_fd_sc_hd__nor2_1 _10424_ (.A(net536),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__mux4_1 _10425_ (.A0(\dpath.RF.R[20][25] ),
    .A1(\dpath.RF.R[21][25] ),
    .A2(\dpath.RF.R[22][25] ),
    .A3(\dpath.RF.R[23][25] ),
    .S0(net570),
    .S1(net551),
    .X(_04618_));
 sky130_fd_sc_hd__nor2_1 _10426_ (.A(net513),
    .B(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__mux4_1 _10427_ (.A0(\dpath.RF.R[28][25] ),
    .A1(\dpath.RF.R[29][25] ),
    .A2(\dpath.RF.R[30][25] ),
    .A3(\dpath.RF.R[31][25] ),
    .S0(net573),
    .S1(net554),
    .X(_04620_));
 sky130_fd_sc_hd__nor2_1 _10428_ (.A(net515),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__mux4_1 _10429_ (.A0(\dpath.RF.R[24][25] ),
    .A1(\dpath.RF.R[25][25] ),
    .A2(\dpath.RF.R[26][25] ),
    .A3(\dpath.RF.R[27][25] ),
    .S0(net569),
    .S1(net550),
    .X(_04622_));
 sky130_fd_sc_hd__o21ai_1 _10430_ (.A1(net534),
    .A2(_04622_),
    .B1(net525),
    .Y(_04623_));
 sky130_fd_sc_hd__o32a_1 _10431_ (.A1(net526),
    .A2(_04617_),
    .A3(_04619_),
    .B1(_04621_),
    .B2(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__a221o_1 _10432_ (.A1(_04610_),
    .A2(_04615_),
    .B1(_04624_),
    .B2(net520),
    .C1(net483),
    .X(_04625_));
 sky130_fd_sc_hd__nor2_1 _10433_ (.A(_02097_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__mux2_2 _10434_ (.A0(net3590),
    .A1(net18),
    .S(net479),
    .X(_04627_));
 sky130_fd_sc_hd__a221o_2 _10435_ (.A1(net667),
    .A2(net369),
    .B1(net368),
    .B2(_04627_),
    .C1(_04626_),
    .X(_04628_));
 sky130_fd_sc_hd__a21oi_1 _10436_ (.A1(_01899_),
    .A2(_04456_),
    .B1(_01894_),
    .Y(_04629_));
 sky130_fd_sc_hd__a31o_1 _10437_ (.A1(_01894_),
    .A2(_01899_),
    .A3(_04456_),
    .B1(net469),
    .X(_04630_));
 sky130_fd_sc_hd__a31o_1 _10438_ (.A1(net789),
    .A2(\dpath.alu.adder.in0[24] ),
    .A3(_04544_),
    .B1(_04543_),
    .X(_04631_));
 sky130_fd_sc_hd__nor2_1 _10439_ (.A(_04569_),
    .B(_04571_),
    .Y(_04632_));
 sky130_fd_sc_hd__a22o_1 _10440_ (.A1(net648),
    .A2(net720),
    .B1(\dpath.alu.adder.in1[25] ),
    .B2(net652),
    .X(_04633_));
 sky130_fd_sc_hd__a21bo_1 _10441_ (.A1(\dpath.alu.adder.in1[25] ),
    .A2(_04465_),
    .B1_N(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__nand2_1 _10442_ (.A(net644),
    .B(net721),
    .Y(_04635_));
 sky130_fd_sc_hd__xor2_1 _10443_ (.A(_04634_),
    .B(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__and2_1 _10444_ (.A(_04466_),
    .B(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__nor2_1 _10445_ (.A(_04466_),
    .B(_04636_),
    .Y(_04638_));
 sky130_fd_sc_hd__or2_1 _10446_ (.A(_04637_),
    .B(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__and4_1 _10447_ (.A(net640),
    .B(net634),
    .C(net723),
    .D(net722),
    .X(_04640_));
 sky130_fd_sc_hd__nand4_1 _10448_ (.A(net640),
    .B(net634),
    .C(net723),
    .D(net722),
    .Y(_04641_));
 sky130_fd_sc_hd__a22o_1 _10449_ (.A1(net634),
    .A2(net723),
    .B1(net722),
    .B2(net640),
    .X(_04642_));
 sky130_fd_sc_hd__and4_1 _10450_ (.A(net630),
    .B(net725),
    .C(_04641_),
    .D(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__a22oi_1 _10451_ (.A1(net630),
    .A2(net725),
    .B1(_04641_),
    .B2(_04642_),
    .Y(_04644_));
 sky130_fd_sc_hd__or2_1 _10452_ (.A(_04643_),
    .B(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__a31o_1 _10453_ (.A1(net634),
    .A2(net725),
    .A3(_04470_),
    .B1(_04469_),
    .X(_04646_));
 sky130_fd_sc_hd__nand2b_1 _10454_ (.A_N(_04645_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__xor2_2 _10455_ (.A(_04645_),
    .B(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__and3_1 _10456_ (.A(net626),
    .B(net622),
    .C(net726),
    .X(_04649_));
 sky130_fd_sc_hd__a22o_1 _10457_ (.A1(net622),
    .A2(net728),
    .B1(net726),
    .B2(net626),
    .X(_04650_));
 sky130_fd_sc_hd__a21bo_1 _10458_ (.A1(net728),
    .A2(_04649_),
    .B1_N(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__nand2_1 _10459_ (.A(net618),
    .B(net730),
    .Y(_04652_));
 sky130_fd_sc_hd__xnor2_1 _10460_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__xor2_1 _10461_ (.A(_04648_),
    .B(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__o21a_1 _10462_ (.A1(_04475_),
    .A2(_04482_),
    .B1(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__nor3_1 _10463_ (.A(_04475_),
    .B(_04482_),
    .C(_04654_),
    .Y(_04656_));
 sky130_fd_sc_hd__or3_2 _10464_ (.A(_04639_),
    .B(_04655_),
    .C(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__o21ai_1 _10465_ (.A1(_04655_),
    .A2(_04656_),
    .B1(_04639_),
    .Y(_04658_));
 sky130_fd_sc_hd__a21o_1 _10466_ (.A1(_04657_),
    .A2(_04658_),
    .B1(_04487_),
    .X(_04659_));
 sky130_fd_sc_hd__nand3_2 _10467_ (.A(_04487_),
    .B(_04657_),
    .C(_04658_),
    .Y(_04660_));
 sky130_fd_sc_hd__and3_1 _10468_ (.A(net756),
    .B(net753),
    .C(net595),
    .X(_04661_));
 sky130_fd_sc_hd__a22o_1 _10469_ (.A1(net753),
    .A2(net596),
    .B1(net592),
    .B2(net756),
    .X(_04662_));
 sky130_fd_sc_hd__a21bo_1 _10470_ (.A1(net592),
    .A2(_04661_),
    .B1_N(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(net759),
    .B(net589),
    .Y(_04664_));
 sky130_fd_sc_hd__xor2_2 _10472_ (.A(_04663_),
    .B(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__and4_1 _10473_ (.A(net604),
    .B(net743),
    .C(net601),
    .D(net739),
    .X(_04666_));
 sky130_fd_sc_hd__nand4_1 _10474_ (.A(net604),
    .B(net743),
    .C(net601),
    .D(net739),
    .Y(_04667_));
 sky130_fd_sc_hd__a22o_1 _10475_ (.A1(net743),
    .A2(net601),
    .B1(net739),
    .B2(net604),
    .X(_04668_));
 sky130_fd_sc_hd__and4_1 _10476_ (.A(net747),
    .B(net598),
    .C(_04667_),
    .D(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__nand4_1 _10477_ (.A(net747),
    .B(net598),
    .C(_04667_),
    .D(_04668_),
    .Y(_04670_));
 sky130_fd_sc_hd__a22o_1 _10478_ (.A1(net747),
    .A2(net598),
    .B1(_04667_),
    .B2(_04668_),
    .X(_04671_));
 sky130_fd_sc_hd__o211a_1 _10479_ (.A1(_04497_),
    .A2(_04499_),
    .B1(_04670_),
    .C1(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__a211o_1 _10480_ (.A1(_04670_),
    .A2(_04671_),
    .B1(_04497_),
    .C1(_04499_),
    .X(_04673_));
 sky130_fd_sc_hd__nand2b_1 _10481_ (.A_N(_04672_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__xnor2_2 _10482_ (.A(_04665_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2_1 _10483_ (.A(_04508_),
    .B(_04510_),
    .Y(_04676_));
 sky130_fd_sc_hd__a21bo_1 _10484_ (.A1(_04478_),
    .A2(_04480_),
    .B1_N(_04477_),
    .X(_04677_));
 sky130_fd_sc_hd__nand4_2 _10485_ (.A(net614),
    .B(net610),
    .C(net735),
    .D(net733),
    .Y(_04678_));
 sky130_fd_sc_hd__a22o_1 _10486_ (.A1(net610),
    .A2(net735),
    .B1(net733),
    .B2(net614),
    .X(_04679_));
 sky130_fd_sc_hd__nand4_2 _10487_ (.A(net609),
    .B(net738),
    .C(_04678_),
    .D(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__a22o_1 _10488_ (.A1(net609),
    .A2(net738),
    .B1(_04678_),
    .B2(_04679_),
    .X(_04681_));
 sky130_fd_sc_hd__nand3_1 _10489_ (.A(_04677_),
    .B(_04680_),
    .C(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__a21o_1 _10490_ (.A1(_04680_),
    .A2(_04681_),
    .B1(_04677_),
    .X(_04683_));
 sky130_fd_sc_hd__nand3_1 _10491_ (.A(_04676_),
    .B(_04682_),
    .C(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__a21o_1 _10492_ (.A1(_04682_),
    .A2(_04683_),
    .B1(_04676_),
    .X(_04685_));
 sky130_fd_sc_hd__a21bo_1 _10493_ (.A1(_04506_),
    .A2(_04513_),
    .B1_N(_04512_),
    .X(_04686_));
 sky130_fd_sc_hd__and3_1 _10494_ (.A(_04684_),
    .B(_04685_),
    .C(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__a21oi_1 _10495_ (.A1(_04684_),
    .A2(_04685_),
    .B1(_04686_),
    .Y(_04688_));
 sky130_fd_sc_hd__nor3b_2 _10496_ (.A(_04687_),
    .B(_04688_),
    .C_N(_04675_),
    .Y(_04689_));
 sky130_fd_sc_hd__o21ba_1 _10497_ (.A1(_04687_),
    .A2(_04688_),
    .B1_N(_04675_),
    .X(_04690_));
 sky130_fd_sc_hd__or3_4 _10498_ (.A(_04485_),
    .B(_04689_),
    .C(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__o21ai_2 _10499_ (.A1(_04689_),
    .A2(_04690_),
    .B1(_04485_),
    .Y(_04692_));
 sky130_fd_sc_hd__o211ai_4 _10500_ (.A1(_04517_),
    .A2(_04520_),
    .B1(_04691_),
    .C1(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__a211o_1 _10501_ (.A1(_04691_),
    .A2(_04692_),
    .B1(_04517_),
    .C1(_04520_),
    .X(_04694_));
 sky130_fd_sc_hd__nand4_4 _10502_ (.A(_04659_),
    .B(_04660_),
    .C(_04693_),
    .D(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__a22o_2 _10503_ (.A1(_04659_),
    .A2(_04660_),
    .B1(_04693_),
    .B2(_04694_),
    .X(_04696_));
 sky130_fd_sc_hd__o211a_1 _10504_ (.A1(_04489_),
    .A2(_04526_),
    .B1(_04695_),
    .C1(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__o211ai_4 _10505_ (.A1(_04489_),
    .A2(_04526_),
    .B1(_04695_),
    .C1(_04696_),
    .Y(_04698_));
 sky130_fd_sc_hd__a211oi_2 _10506_ (.A1(_04695_),
    .A2(_04696_),
    .B1(_04489_),
    .C1(_04526_),
    .Y(_04699_));
 sky130_fd_sc_hd__nand4_2 _10507_ (.A(net776),
    .B(net775),
    .C(net581),
    .D(net580),
    .Y(_04700_));
 sky130_fd_sc_hd__a22o_1 _10508_ (.A1(net772),
    .A2(net581),
    .B1(net580),
    .B2(net776),
    .X(_04701_));
 sky130_fd_sc_hd__and2_1 _10509_ (.A(net780),
    .B(net579),
    .X(_04702_));
 sky130_fd_sc_hd__nand3_1 _10510_ (.A(_04700_),
    .B(_04701_),
    .C(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__a21o_1 _10511_ (.A1(_04700_),
    .A2(_04701_),
    .B1(_04702_),
    .X(_04704_));
 sky130_fd_sc_hd__a31o_1 _10512_ (.A1(net782),
    .A2(net580),
    .A3(_04533_),
    .B1(_04532_),
    .X(_04705_));
 sky130_fd_sc_hd__and3_1 _10513_ (.A(_04703_),
    .B(_04704_),
    .C(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__a21oi_1 _10514_ (.A1(_04703_),
    .A2(_04704_),
    .B1(_04705_),
    .Y(_04707_));
 sky130_fd_sc_hd__or2_1 _10515_ (.A(_04706_),
    .B(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__nand2_1 _10516_ (.A(net784),
    .B(\dpath.alu.adder.in0[24] ),
    .Y(_04709_));
 sky130_fd_sc_hd__xor2_2 _10517_ (.A(_04708_),
    .B(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__a31o_1 _10518_ (.A1(net784),
    .A2(\dpath.alu.adder.in0[23] ),
    .A3(_04539_),
    .B1(_04538_),
    .X(_04711_));
 sky130_fd_sc_hd__xor2_2 _10519_ (.A(_04710_),
    .B(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__nand2_1 _10520_ (.A(net787),
    .B(\dpath.alu.adder.in0[25] ),
    .Y(_04713_));
 sky130_fd_sc_hd__and3_1 _10521_ (.A(net787),
    .B(\dpath.alu.adder.in0[25] ),
    .C(_04712_),
    .X(_04714_));
 sky130_fd_sc_hd__xor2_2 _10522_ (.A(_04712_),
    .B(_04713_),
    .X(_04715_));
 sky130_fd_sc_hd__a21o_1 _10523_ (.A1(_04495_),
    .A2(_04503_),
    .B1(_04502_),
    .X(_04716_));
 sky130_fd_sc_hd__nand2_1 _10524_ (.A(_04550_),
    .B(_04552_),
    .Y(_04717_));
 sky130_fd_sc_hd__a32o_1 _10525_ (.A1(net759),
    .A2(net592),
    .A3(_04492_),
    .B1(_04491_),
    .B2(net595),
    .X(_04718_));
 sky130_fd_sc_hd__nand4_2 _10526_ (.A(net764),
    .B(net760),
    .C(net587),
    .D(net585),
    .Y(_04719_));
 sky130_fd_sc_hd__a22o_1 _10527_ (.A1(net763),
    .A2(net587),
    .B1(net585),
    .B2(\dpath.alu.adder.in1[6] ),
    .X(_04720_));
 sky130_fd_sc_hd__nand4_2 _10528_ (.A(net768),
    .B(net583),
    .C(_04719_),
    .D(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__a22o_1 _10529_ (.A1(net768),
    .A2(net583),
    .B1(_04719_),
    .B2(_04720_),
    .X(_04722_));
 sky130_fd_sc_hd__nand3_2 _10530_ (.A(_04718_),
    .B(_04721_),
    .C(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__a21o_1 _10531_ (.A1(_04721_),
    .A2(_04722_),
    .B1(_04718_),
    .X(_04724_));
 sky130_fd_sc_hd__nand3_2 _10532_ (.A(_04717_),
    .B(_04723_),
    .C(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__a21o_1 _10533_ (.A1(_04723_),
    .A2(_04724_),
    .B1(_04717_),
    .X(_04726_));
 sky130_fd_sc_hd__and3_2 _10534_ (.A(_04716_),
    .B(_04725_),
    .C(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__a21oi_2 _10535_ (.A1(_04725_),
    .A2(_04726_),
    .B1(_04716_),
    .Y(_04728_));
 sky130_fd_sc_hd__a211oi_1 _10536_ (.A1(_04554_),
    .A2(_04556_),
    .B1(_04727_),
    .C1(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__a211o_1 _10537_ (.A1(_04554_),
    .A2(_04556_),
    .B1(_04727_),
    .C1(_04728_),
    .X(_04730_));
 sky130_fd_sc_hd__o211ai_2 _10538_ (.A1(_04727_),
    .A2(_04728_),
    .B1(_04554_),
    .C1(_04556_),
    .Y(_04731_));
 sky130_fd_sc_hd__o211a_1 _10539_ (.A1(_04558_),
    .A2(_04560_),
    .B1(_04730_),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__a211oi_2 _10540_ (.A1(_04730_),
    .A2(_04731_),
    .B1(_04558_),
    .C1(_04560_),
    .Y(_04733_));
 sky130_fd_sc_hd__nor3_2 _10541_ (.A(_04715_),
    .B(_04732_),
    .C(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__o21a_1 _10542_ (.A1(_04732_),
    .A2(_04733_),
    .B1(_04715_),
    .X(_04735_));
 sky130_fd_sc_hd__a211oi_4 _10543_ (.A1(_04522_),
    .A2(_04524_),
    .B1(_04734_),
    .C1(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__o211a_1 _10544_ (.A1(_04734_),
    .A2(_04735_),
    .B1(_04522_),
    .C1(_04524_),
    .X(_04737_));
 sky130_fd_sc_hd__a211oi_4 _10545_ (.A1(_04564_),
    .A2(_04567_),
    .B1(_04736_),
    .C1(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__o211a_1 _10546_ (.A1(_04736_),
    .A2(_04737_),
    .B1(_04564_),
    .C1(_04567_),
    .X(_04739_));
 sky130_fd_sc_hd__nor4_1 _10547_ (.A(_04697_),
    .B(_04699_),
    .C(_04738_),
    .D(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__or4_2 _10548_ (.A(_04697_),
    .B(_04699_),
    .C(_04738_),
    .D(_04739_),
    .X(_04741_));
 sky130_fd_sc_hd__o22a_1 _10549_ (.A1(_04697_),
    .A2(_04699_),
    .B1(_04738_),
    .B2(_04739_),
    .X(_04742_));
 sky130_fd_sc_hd__a211oi_2 _10550_ (.A1(_04531_),
    .A2(_04574_),
    .B1(_04740_),
    .C1(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__o211a_1 _10551_ (.A1(_04740_),
    .A2(_04742_),
    .B1(_04531_),
    .C1(_04574_),
    .X(_04744_));
 sky130_fd_sc_hd__nor3_1 _10552_ (.A(_04632_),
    .B(_04743_),
    .C(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__or3_1 _10553_ (.A(_04632_),
    .B(_04743_),
    .C(_04744_),
    .X(_04746_));
 sky130_fd_sc_hd__o21ai_1 _10554_ (.A1(_04743_),
    .A2(_04744_),
    .B1(_04632_),
    .Y(_04747_));
 sky130_fd_sc_hd__o211a_1 _10555_ (.A1(_04576_),
    .A2(_04578_),
    .B1(_04746_),
    .C1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__a211oi_1 _10556_ (.A1(_04746_),
    .A2(_04747_),
    .B1(_04576_),
    .C1(_04578_),
    .Y(_04749_));
 sky130_fd_sc_hd__nor2_1 _10557_ (.A(_04748_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__xor2_1 _10558_ (.A(_04631_),
    .B(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__o21a_1 _10559_ (.A1(_04581_),
    .A2(_04583_),
    .B1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__or3_1 _10560_ (.A(_04581_),
    .B(_04583_),
    .C(_04751_),
    .X(_04753_));
 sky130_fd_sc_hd__and2b_1 _10561_ (.A_N(_04752_),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__nor2_1 _10562_ (.A(_04587_),
    .B(_04590_),
    .Y(_04755_));
 sky130_fd_sc_hd__xor2_1 _10563_ (.A(_04754_),
    .B(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__nor2_1 _10564_ (.A(net3691),
    .B(_02071_),
    .Y(_04757_));
 sky130_fd_sc_hd__a211o_1 _10565_ (.A1(net484),
    .A2(_04756_),
    .B1(_04757_),
    .C1(net467),
    .X(_04758_));
 sky130_fd_sc_hd__o21ai_4 _10566_ (.A1(_04629_),
    .A2(_04630_),
    .B1(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__a21oi_4 _10567_ (.A1(net391),
    .A2(_04759_),
    .B1(_04628_),
    .Y(_04760_));
 sky130_fd_sc_hd__xnor2_1 _10568_ (.A(net577),
    .B(net3522),
    .Y(_04761_));
 sky130_fd_sc_hd__o21a_1 _10569_ (.A1(_04597_),
    .A2(_04600_),
    .B1(_04599_),
    .X(_04762_));
 sky130_fd_sc_hd__xnor2_1 _10570_ (.A(_04761_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_1 _10571_ (.A(_01760_),
    .B(_04603_),
    .Y(_04764_));
 sky130_fd_sc_hd__a211o_1 _10572_ (.A1(_01760_),
    .A2(_04603_),
    .B1(_04764_),
    .C1(_01958_),
    .X(_04765_));
 sky130_fd_sc_hd__a21oi_1 _10573_ (.A1(\dpath.btarg_DX.q[25] ),
    .A2(net404),
    .B1(net451),
    .Y(_04766_));
 sky130_fd_sc_hd__o211a_1 _10574_ (.A1(net366),
    .A2(_04763_),
    .B1(_04765_),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__o21ai_1 _10575_ (.A1(net374),
    .A2(_04760_),
    .B1(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__o211a_1 _10576_ (.A1(net3507),
    .A2(net443),
    .B1(_04768_),
    .C1(net852),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_1 _10577_ (.A0(\dpath.RF.R[0][26] ),
    .A1(\dpath.RF.R[1][26] ),
    .A2(\dpath.RF.R[2][26] ),
    .A3(\dpath.RF.R[3][26] ),
    .S0(net571),
    .S1(net552),
    .X(_04769_));
 sky130_fd_sc_hd__mux4_1 _10578_ (.A0(\dpath.RF.R[4][26] ),
    .A1(\dpath.RF.R[5][26] ),
    .A2(\dpath.RF.R[6][26] ),
    .A3(\dpath.RF.R[7][26] ),
    .S0(net571),
    .S1(net552),
    .X(_04770_));
 sky130_fd_sc_hd__o21a_1 _10579_ (.A1(net516),
    .A2(_04770_),
    .B1(net507),
    .X(_04771_));
 sky130_fd_sc_hd__o21ai_1 _10580_ (.A1(net537),
    .A2(_04769_),
    .B1(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__mux4_1 _10581_ (.A0(\dpath.RF.R[12][26] ),
    .A1(\dpath.RF.R[13][26] ),
    .A2(\dpath.RF.R[14][26] ),
    .A3(\dpath.RF.R[15][26] ),
    .S0(net571),
    .S1(net552),
    .X(_04773_));
 sky130_fd_sc_hd__mux4_1 _10582_ (.A0(\dpath.RF.R[8][26] ),
    .A1(\dpath.RF.R[9][26] ),
    .A2(\dpath.RF.R[10][26] ),
    .A3(\dpath.RF.R[11][26] ),
    .S0(net571),
    .S1(net552),
    .X(_04774_));
 sky130_fd_sc_hd__or2_1 _10583_ (.A(net537),
    .B(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__o211a_1 _10584_ (.A1(net516),
    .A2(_04773_),
    .B1(_04775_),
    .C1(net527),
    .X(_04776_));
 sky130_fd_sc_hd__nor2_1 _10585_ (.A(net520),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__mux4_1 _10586_ (.A0(\dpath.RF.R[16][26] ),
    .A1(\dpath.RF.R[17][26] ),
    .A2(\dpath.RF.R[18][26] ),
    .A3(\dpath.RF.R[19][26] ),
    .S0(net572),
    .S1(net553),
    .X(_04778_));
 sky130_fd_sc_hd__nor2_1 _10587_ (.A(net537),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__mux4_1 _10588_ (.A0(\dpath.RF.R[20][26] ),
    .A1(\dpath.RF.R[21][26] ),
    .A2(\dpath.RF.R[22][26] ),
    .A3(\dpath.RF.R[23][26] ),
    .S0(net572),
    .S1(net553),
    .X(_04780_));
 sky130_fd_sc_hd__nor2_1 _10589_ (.A(net516),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__mux4_1 _10590_ (.A0(\dpath.RF.R[28][26] ),
    .A1(\dpath.RF.R[29][26] ),
    .A2(\dpath.RF.R[30][26] ),
    .A3(\dpath.RF.R[31][26] ),
    .S0(net572),
    .S1(net553),
    .X(_04782_));
 sky130_fd_sc_hd__nor2_1 _10591_ (.A(net516),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__mux4_1 _10592_ (.A0(\dpath.RF.R[24][26] ),
    .A1(\dpath.RF.R[25][26] ),
    .A2(\dpath.RF.R[26][26] ),
    .A3(\dpath.RF.R[27][26] ),
    .S0(net572),
    .S1(net553),
    .X(_04784_));
 sky130_fd_sc_hd__o21ai_1 _10593_ (.A1(net537),
    .A2(_04784_),
    .B1(net527),
    .Y(_04785_));
 sky130_fd_sc_hd__o32a_1 _10594_ (.A1(net527),
    .A2(_04779_),
    .A3(_04781_),
    .B1(_04783_),
    .B2(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__a221o_1 _10595_ (.A1(_04772_),
    .A2(_04777_),
    .B1(_04786_),
    .B2(net520),
    .C1(net483),
    .X(_04787_));
 sky130_fd_sc_hd__nor2_1 _10596_ (.A(net371),
    .B(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__mux2_2 _10597_ (.A0(net3655),
    .A1(net19),
    .S(net480),
    .X(_04789_));
 sky130_fd_sc_hd__a221o_1 _10598_ (.A1(net664),
    .A2(net369),
    .B1(net367),
    .B2(_04789_),
    .C1(_04788_),
    .X(_04790_));
 sky130_fd_sc_hd__a21bo_1 _10599_ (.A1(_01893_),
    .A2(_01899_),
    .B1_N(_01892_),
    .X(_04791_));
 sky130_fd_sc_hd__or2_1 _10600_ (.A(_01894_),
    .B(_01900_),
    .X(_04792_));
 sky130_fd_sc_hd__or2_1 _10601_ (.A(_04454_),
    .B(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__a21o_1 _10602_ (.A1(_04791_),
    .A2(_04793_),
    .B1(_01916_),
    .X(_04794_));
 sky130_fd_sc_hd__a21oi_1 _10603_ (.A1(_04710_),
    .A2(_04711_),
    .B1(_04714_),
    .Y(_04795_));
 sky130_fd_sc_hd__nand2_1 _10604_ (.A(net652),
    .B(\dpath.alu.adder.in1[26] ),
    .Y(_04796_));
 sky130_fd_sc_hd__a22oi_1 _10605_ (.A1(net644),
    .A2(net720),
    .B1(\dpath.alu.adder.in1[25] ),
    .B2(net648),
    .Y(_04797_));
 sky130_fd_sc_hd__and4_1 _10606_ (.A(net648),
    .B(net644),
    .C(net720),
    .D(\dpath.alu.adder.in1[25] ),
    .X(_04798_));
 sky130_fd_sc_hd__o2bb2a_1 _10607_ (.A1_N(net640),
    .A2_N(net721),
    .B1(_04797_),
    .B2(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__and4bb_1 _10608_ (.A_N(_04797_),
    .B_N(_04798_),
    .C(net640),
    .D(net721),
    .X(_04800_));
 sky130_fd_sc_hd__or2_1 _10609_ (.A(_04799_),
    .B(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__a32o_1 _10610_ (.A1(net644),
    .A2(net721),
    .A3(_04633_),
    .B1(_04465_),
    .B2(\dpath.alu.adder.in1[25] ),
    .X(_04802_));
 sky130_fd_sc_hd__and2b_1 _10611_ (.A_N(_04801_),
    .B(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__xnor2_1 _10612_ (.A(_04801_),
    .B(_04802_),
    .Y(_04804_));
 sky130_fd_sc_hd__nand2b_1 _10613_ (.A_N(_04796_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__xnor2_1 _10614_ (.A(_04796_),
    .B(_04804_),
    .Y(_04806_));
 sky130_fd_sc_hd__o21ai_2 _10615_ (.A1(_04648_),
    .A2(_04653_),
    .B1(_04647_),
    .Y(_04807_));
 sky130_fd_sc_hd__a22o_1 _10616_ (.A1(net618),
    .A2(net728),
    .B1(net726),
    .B2(net622),
    .X(_04808_));
 sky130_fd_sc_hd__nand4_4 _10617_ (.A(net622),
    .B(net618),
    .C(net728),
    .D(net726),
    .Y(_04809_));
 sky130_fd_sc_hd__a22o_1 _10618_ (.A1(net614),
    .A2(net730),
    .B1(_04808_),
    .B2(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__nand4_2 _10619_ (.A(net614),
    .B(net730),
    .C(_04808_),
    .D(_04809_),
    .Y(_04811_));
 sky130_fd_sc_hd__and2_1 _10620_ (.A(_04810_),
    .B(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__nand4_4 _10621_ (.A(net634),
    .B(net630),
    .C(net723),
    .D(net722),
    .Y(_04813_));
 sky130_fd_sc_hd__a22o_1 _10622_ (.A1(net630),
    .A2(net723),
    .B1(net722),
    .B2(net634),
    .X(_04814_));
 sky130_fd_sc_hd__nand4_4 _10623_ (.A(net626),
    .B(net725),
    .C(_04813_),
    .D(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__a22o_1 _10624_ (.A1(net626),
    .A2(net725),
    .B1(_04813_),
    .B2(_04814_),
    .X(_04816_));
 sky130_fd_sc_hd__o211ai_4 _10625_ (.A1(_04640_),
    .A2(_04643_),
    .B1(_04815_),
    .C1(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__a211o_1 _10626_ (.A1(_04815_),
    .A2(_04816_),
    .B1(_04640_),
    .C1(_04643_),
    .X(_04818_));
 sky130_fd_sc_hd__nand3_2 _10627_ (.A(_04812_),
    .B(_04817_),
    .C(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__a21o_1 _10628_ (.A1(_04817_),
    .A2(_04818_),
    .B1(_04812_),
    .X(_04820_));
 sky130_fd_sc_hd__nand3_4 _10629_ (.A(_04637_),
    .B(_04819_),
    .C(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21o_1 _10630_ (.A1(_04819_),
    .A2(_04820_),
    .B1(_04637_),
    .X(_04822_));
 sky130_fd_sc_hd__nand3_2 _10631_ (.A(_04807_),
    .B(_04821_),
    .C(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__a21o_1 _10632_ (.A1(_04821_),
    .A2(_04822_),
    .B1(_04807_),
    .X(_04824_));
 sky130_fd_sc_hd__and3_1 _10633_ (.A(_04806_),
    .B(_04823_),
    .C(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__a21oi_1 _10634_ (.A1(_04823_),
    .A2(_04824_),
    .B1(_04806_),
    .Y(_04826_));
 sky130_fd_sc_hd__nor3_2 _10635_ (.A(_04657_),
    .B(_04825_),
    .C(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__o21a_1 _10636_ (.A1(_04825_),
    .A2(_04826_),
    .B1(_04657_),
    .X(_04828_));
 sky130_fd_sc_hd__nand4_4 _10637_ (.A(net756),
    .B(net753),
    .C(net593),
    .D(net589),
    .Y(_04829_));
 sky130_fd_sc_hd__a22o_1 _10638_ (.A1(net753),
    .A2(net593),
    .B1(net589),
    .B2(net756),
    .X(_04830_));
 sky130_fd_sc_hd__nand4_2 _10639_ (.A(net759),
    .B(net587),
    .C(_04829_),
    .D(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__a22o_1 _10640_ (.A1(net759),
    .A2(net587),
    .B1(_04829_),
    .B2(_04830_),
    .X(_04832_));
 sky130_fd_sc_hd__and2_1 _10641_ (.A(_04831_),
    .B(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__and4_1 _10642_ (.A(net743),
    .B(net601),
    .C(\dpath.alu.adder.in1[13] ),
    .D(net598),
    .X(_04834_));
 sky130_fd_sc_hd__nand4_2 _10643_ (.A(net743),
    .B(net601),
    .C(net739),
    .D(net598),
    .Y(_04835_));
 sky130_fd_sc_hd__a22o_1 _10644_ (.A1(net601),
    .A2(net739),
    .B1(net598),
    .B2(net743),
    .X(_04836_));
 sky130_fd_sc_hd__and4_1 _10645_ (.A(net747),
    .B(net595),
    .C(_04835_),
    .D(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__nand4_1 _10646_ (.A(net747),
    .B(net595),
    .C(_04835_),
    .D(_04836_),
    .Y(_04838_));
 sky130_fd_sc_hd__a22o_1 _10647_ (.A1(net747),
    .A2(net596),
    .B1(_04835_),
    .B2(_04836_),
    .X(_04839_));
 sky130_fd_sc_hd__o211a_1 _10648_ (.A1(_04666_),
    .A2(_04669_),
    .B1(_04838_),
    .C1(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__a211o_1 _10649_ (.A1(_04838_),
    .A2(_04839_),
    .B1(_04666_),
    .C1(_04669_),
    .X(_04841_));
 sky130_fd_sc_hd__nand2b_1 _10650_ (.A_N(_04840_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__xnor2_2 _10651_ (.A(_04833_),
    .B(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_1 _10652_ (.A(_04678_),
    .B(_04680_),
    .Y(_04844_));
 sky130_fd_sc_hd__a32o_1 _10653_ (.A1(net618),
    .A2(net730),
    .A3(_04650_),
    .B1(_04649_),
    .B2(net729),
    .X(_04845_));
 sky130_fd_sc_hd__nand4_1 _10654_ (.A(net610),
    .B(net607),
    .C(net735),
    .D(net733),
    .Y(_04846_));
 sky130_fd_sc_hd__a22o_1 _10655_ (.A1(net607),
    .A2(net735),
    .B1(net733),
    .B2(\dpath.alu.adder.in0[10] ),
    .X(_04847_));
 sky130_fd_sc_hd__nand4_1 _10656_ (.A(net605),
    .B(net738),
    .C(_04846_),
    .D(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__a22o_1 _10657_ (.A1(net605),
    .A2(net738),
    .B1(_04846_),
    .B2(_04847_),
    .X(_04849_));
 sky130_fd_sc_hd__nand3_1 _10658_ (.A(_04845_),
    .B(_04848_),
    .C(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__a21o_1 _10659_ (.A1(_04848_),
    .A2(_04849_),
    .B1(_04845_),
    .X(_04851_));
 sky130_fd_sc_hd__nand3_1 _10660_ (.A(_04844_),
    .B(_04850_),
    .C(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__a21o_1 _10661_ (.A1(_04850_),
    .A2(_04851_),
    .B1(_04844_),
    .X(_04853_));
 sky130_fd_sc_hd__a21bo_1 _10662_ (.A1(_04676_),
    .A2(_04683_),
    .B1_N(_04682_),
    .X(_04854_));
 sky130_fd_sc_hd__and3_1 _10663_ (.A(_04852_),
    .B(_04853_),
    .C(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__nand3_1 _10664_ (.A(_04852_),
    .B(_04853_),
    .C(_04854_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21o_1 _10665_ (.A1(_04852_),
    .A2(_04853_),
    .B1(_04854_),
    .X(_04857_));
 sky130_fd_sc_hd__and3_2 _10666_ (.A(_04843_),
    .B(_04856_),
    .C(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__a21oi_1 _10667_ (.A1(_04856_),
    .A2(_04857_),
    .B1(_04843_),
    .Y(_04859_));
 sky130_fd_sc_hd__or3b_2 _10668_ (.A(_04858_),
    .B(_04859_),
    .C_N(_04655_),
    .X(_04860_));
 sky130_fd_sc_hd__inv_2 _10669_ (.A(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__o21bai_1 _10670_ (.A1(_04858_),
    .A2(_04859_),
    .B1_N(_04655_),
    .Y(_04862_));
 sky130_fd_sc_hd__o211a_1 _10671_ (.A1(_04687_),
    .A2(_04689_),
    .B1(_04860_),
    .C1(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__a211oi_1 _10672_ (.A1(_04860_),
    .A2(_04862_),
    .B1(_04687_),
    .C1(_04689_),
    .Y(_04864_));
 sky130_fd_sc_hd__nor4_2 _10673_ (.A(_04827_),
    .B(_04828_),
    .C(_04863_),
    .D(_04864_),
    .Y(_04865_));
 sky130_fd_sc_hd__o22a_1 _10674_ (.A1(_04827_),
    .A2(_04828_),
    .B1(_04863_),
    .B2(_04864_),
    .X(_04866_));
 sky130_fd_sc_hd__a211oi_2 _10675_ (.A1(_04660_),
    .A2(_04695_),
    .B1(_04865_),
    .C1(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__o211a_1 _10676_ (.A1(_04865_),
    .A2(_04866_),
    .B1(_04660_),
    .C1(_04695_),
    .X(_04868_));
 sky130_fd_sc_hd__or2_1 _10677_ (.A(_04732_),
    .B(_04734_),
    .X(_04869_));
 sky130_fd_sc_hd__nand4_1 _10678_ (.A(net777),
    .B(net772),
    .C(\dpath.alu.adder.in0[22] ),
    .D(net579),
    .Y(_04870_));
 sky130_fd_sc_hd__a22o_1 _10679_ (.A1(net772),
    .A2(\dpath.alu.adder.in0[22] ),
    .B1(net579),
    .B2(net777),
    .X(_04871_));
 sky130_fd_sc_hd__and2_1 _10680_ (.A(net780),
    .B(\dpath.alu.adder.in0[24] ),
    .X(_04872_));
 sky130_fd_sc_hd__nand3_1 _10681_ (.A(_04870_),
    .B(_04871_),
    .C(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__a21o_1 _10682_ (.A1(_04870_),
    .A2(_04871_),
    .B1(_04872_),
    .X(_04874_));
 sky130_fd_sc_hd__a21bo_1 _10683_ (.A1(_04701_),
    .A2(_04702_),
    .B1_N(_04700_),
    .X(_04875_));
 sky130_fd_sc_hd__and3_1 _10684_ (.A(_04873_),
    .B(_04874_),
    .C(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__a21oi_1 _10685_ (.A1(_04873_),
    .A2(_04874_),
    .B1(_04875_),
    .Y(_04877_));
 sky130_fd_sc_hd__or2_1 _10686_ (.A(_04876_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _10687_ (.A(net784),
    .B(\dpath.alu.adder.in0[25] ),
    .Y(_04879_));
 sky130_fd_sc_hd__xnor2_1 _10688_ (.A(_04878_),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__o21ba_1 _10689_ (.A1(_04707_),
    .A2(_04709_),
    .B1_N(_04706_),
    .X(_04881_));
 sky130_fd_sc_hd__or2_1 _10690_ (.A(_04880_),
    .B(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__xor2_1 _10691_ (.A(_04880_),
    .B(_04881_),
    .X(_04883_));
 sky130_fd_sc_hd__nand2_1 _10692_ (.A(net787),
    .B(\dpath.alu.adder.in0[26] ),
    .Y(_04884_));
 sky130_fd_sc_hd__nand3_1 _10693_ (.A(net786),
    .B(\dpath.alu.adder.in0[26] ),
    .C(_04883_),
    .Y(_04885_));
 sky130_fd_sc_hd__xor2_1 _10694_ (.A(_04883_),
    .B(_04884_),
    .X(_04886_));
 sky130_fd_sc_hd__a21o_1 _10695_ (.A1(_04665_),
    .A2(_04673_),
    .B1(_04672_),
    .X(_04887_));
 sky130_fd_sc_hd__nand2_1 _10696_ (.A(_04719_),
    .B(_04721_),
    .Y(_04888_));
 sky130_fd_sc_hd__a32o_1 _10697_ (.A1(net759),
    .A2(net589),
    .A3(_04662_),
    .B1(_04661_),
    .B2(net592),
    .X(_04889_));
 sky130_fd_sc_hd__nand4_2 _10698_ (.A(\dpath.alu.adder.in1[6] ),
    .B(net763),
    .C(net585),
    .D(net583),
    .Y(_04890_));
 sky130_fd_sc_hd__a22o_1 _10699_ (.A1(net763),
    .A2(net585),
    .B1(net583),
    .B2(\dpath.alu.adder.in1[6] ),
    .X(_04891_));
 sky130_fd_sc_hd__nand4_2 _10700_ (.A(net771),
    .B(net581),
    .C(_04890_),
    .D(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__a22o_1 _10701_ (.A1(net771),
    .A2(net581),
    .B1(_04890_),
    .B2(_04891_),
    .X(_04893_));
 sky130_fd_sc_hd__nand3_2 _10702_ (.A(_04889_),
    .B(_04892_),
    .C(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__a21o_1 _10703_ (.A1(_04892_),
    .A2(_04893_),
    .B1(_04889_),
    .X(_04895_));
 sky130_fd_sc_hd__nand3_2 _10704_ (.A(_04888_),
    .B(_04894_),
    .C(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__a21o_1 _10705_ (.A1(_04894_),
    .A2(_04895_),
    .B1(_04888_),
    .X(_04897_));
 sky130_fd_sc_hd__and3_1 _10706_ (.A(_04887_),
    .B(_04896_),
    .C(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__nand3_1 _10707_ (.A(_04887_),
    .B(_04896_),
    .C(_04897_),
    .Y(_04899_));
 sky130_fd_sc_hd__a21oi_1 _10708_ (.A1(_04896_),
    .A2(_04897_),
    .B1(_04887_),
    .Y(_04900_));
 sky130_fd_sc_hd__a211o_1 _10709_ (.A1(_04723_),
    .A2(_04725_),
    .B1(_04898_),
    .C1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__o211ai_2 _10710_ (.A1(_04898_),
    .A2(_04900_),
    .B1(_04723_),
    .C1(_04725_),
    .Y(_04902_));
 sky130_fd_sc_hd__o211a_2 _10711_ (.A1(_04727_),
    .A2(_04729_),
    .B1(_04901_),
    .C1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__a211oi_2 _10712_ (.A1(_04901_),
    .A2(_04902_),
    .B1(_04727_),
    .C1(_04729_),
    .Y(_04904_));
 sky130_fd_sc_hd__nor3_2 _10713_ (.A(_04886_),
    .B(_04903_),
    .C(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__o21a_1 _10714_ (.A1(_04903_),
    .A2(_04904_),
    .B1(_04886_),
    .X(_04906_));
 sky130_fd_sc_hd__a211o_1 _10715_ (.A1(_04691_),
    .A2(_04693_),
    .B1(_04905_),
    .C1(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__o211ai_2 _10716_ (.A1(_04905_),
    .A2(_04906_),
    .B1(_04691_),
    .C1(_04693_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand3_2 _10717_ (.A(_04869_),
    .B(_04907_),
    .C(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__a21o_1 _10718_ (.A1(_04907_),
    .A2(_04908_),
    .B1(_04869_),
    .X(_04910_));
 sky130_fd_sc_hd__and4bb_2 _10719_ (.A_N(_04867_),
    .B_N(_04868_),
    .C(_04909_),
    .D(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__a2bb2oi_2 _10720_ (.A1_N(_04867_),
    .A2_N(_04868_),
    .B1(_04909_),
    .B2(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__a211o_2 _10721_ (.A1(_04698_),
    .A2(_04741_),
    .B1(_04911_),
    .C1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__o211ai_4 _10722_ (.A1(_04911_),
    .A2(_04912_),
    .B1(_04698_),
    .C1(_04741_),
    .Y(_04914_));
 sky130_fd_sc_hd__o211ai_4 _10723_ (.A1(_04736_),
    .A2(_04738_),
    .B1(_04913_),
    .C1(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__a211o_1 _10724_ (.A1(_04913_),
    .A2(_04914_),
    .B1(_04736_),
    .C1(_04738_),
    .X(_04916_));
 sky130_fd_sc_hd__o211a_1 _10725_ (.A1(_04743_),
    .A2(_04745_),
    .B1(_04915_),
    .C1(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__inv_2 _10726_ (.A(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__a211oi_1 _10727_ (.A1(_04915_),
    .A2(_04916_),
    .B1(_04743_),
    .C1(_04745_),
    .Y(_04919_));
 sky130_fd_sc_hd__or3_1 _10728_ (.A(_04795_),
    .B(_04917_),
    .C(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__o21ai_1 _10729_ (.A1(_04917_),
    .A2(_04919_),
    .B1(_04795_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_1 _10730_ (.A(_04920_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__a21oi_1 _10731_ (.A1(_04631_),
    .A2(_04750_),
    .B1(_04748_),
    .Y(_04923_));
 sky130_fd_sc_hd__or2_1 _10732_ (.A(_04922_),
    .B(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__nand2_1 _10733_ (.A(_04922_),
    .B(_04923_),
    .Y(_04925_));
 sky130_fd_sc_hd__nand2_1 _10734_ (.A(_04924_),
    .B(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__o21ai_1 _10735_ (.A1(_04587_),
    .A2(_04752_),
    .B1(_04753_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2_1 _10736_ (.A(_04588_),
    .B(_04754_),
    .Y(_04928_));
 sky130_fd_sc_hd__o21a_1 _10737_ (.A1(_04462_),
    .A2(_04928_),
    .B1(_04927_),
    .X(_04929_));
 sky130_fd_sc_hd__o21ai_1 _10738_ (.A1(_04926_),
    .A2(_04929_),
    .B1(_02239_),
    .Y(_04930_));
 sky130_fd_sc_hd__a21oi_1 _10739_ (.A1(_04926_),
    .A2(_04929_),
    .B1(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__a31oi_1 _10740_ (.A1(_01916_),
    .A2(_04791_),
    .A3(_04793_),
    .B1(net469),
    .Y(_04932_));
 sky130_fd_sc_hd__a221o_2 _10741_ (.A1(net3601),
    .A2(net486),
    .B1(_04794_),
    .B2(_04932_),
    .C1(_04931_),
    .X(_04933_));
 sky130_fd_sc_hd__a21o_2 _10742_ (.A1(net391),
    .A2(_04933_),
    .B1(_04790_),
    .X(_04934_));
 sky130_fd_sc_hd__or2_1 _10743_ (.A(net577),
    .B(net3509),
    .X(_04935_));
 sky130_fd_sc_hd__nand2_1 _10744_ (.A(net577),
    .B(net3509),
    .Y(_04936_));
 sky130_fd_sc_hd__nand2_1 _10745_ (.A(_04935_),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__or2_1 _10746_ (.A(_04600_),
    .B(_04761_),
    .X(_04938_));
 sky130_fd_sc_hd__o21a_1 _10747_ (.A1(net3522),
    .A2(net3542),
    .B1(net577),
    .X(_04939_));
 sky130_fd_sc_hd__o21ba_1 _10748_ (.A1(_04597_),
    .A2(_04938_),
    .B1_N(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__xnor2_1 _10749_ (.A(_04937_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__nor2_1 _10750_ (.A(net366),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__and2_1 _10751_ (.A(net3368),
    .B(_04764_),
    .X(_04943_));
 sky130_fd_sc_hd__inv_2 _10752_ (.A(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__o211a_1 _10753_ (.A1(net3368),
    .A2(_04764_),
    .B1(_04944_),
    .C1(net362),
    .X(_04945_));
 sky130_fd_sc_hd__a211o_1 _10754_ (.A1(\dpath.btarg_DX.q[26] ),
    .A2(net404),
    .B1(net451),
    .C1(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__a211o_1 _10755_ (.A1(_02027_),
    .A2(_04934_),
    .B1(_04942_),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__o211a_1 _10756_ (.A1(net3368),
    .A2(net444),
    .B1(_04947_),
    .C1(net852),
    .X(_00662_));
 sky130_fd_sc_hd__mux4_1 _10757_ (.A0(\dpath.RF.R[0][27] ),
    .A1(\dpath.RF.R[1][27] ),
    .A2(\dpath.RF.R[2][27] ),
    .A3(\dpath.RF.R[3][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04948_));
 sky130_fd_sc_hd__mux4_1 _10758_ (.A0(\dpath.RF.R[4][27] ),
    .A1(\dpath.RF.R[5][27] ),
    .A2(\dpath.RF.R[6][27] ),
    .A3(\dpath.RF.R[7][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04949_));
 sky130_fd_sc_hd__o21a_1 _10759_ (.A1(net515),
    .A2(_04949_),
    .B1(net507),
    .X(_04950_));
 sky130_fd_sc_hd__o21ai_1 _10760_ (.A1(net536),
    .A2(_04948_),
    .B1(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__mux4_1 _10761_ (.A0(\dpath.RF.R[12][27] ),
    .A1(\dpath.RF.R[13][27] ),
    .A2(\dpath.RF.R[14][27] ),
    .A3(\dpath.RF.R[15][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04952_));
 sky130_fd_sc_hd__mux4_1 _10762_ (.A0(\dpath.RF.R[8][27] ),
    .A1(\dpath.RF.R[9][27] ),
    .A2(\dpath.RF.R[10][27] ),
    .A3(\dpath.RF.R[11][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04953_));
 sky130_fd_sc_hd__or2_1 _10763_ (.A(net536),
    .B(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__o211a_1 _10764_ (.A1(net515),
    .A2(_04952_),
    .B1(_04954_),
    .C1(net526),
    .X(_04955_));
 sky130_fd_sc_hd__nor2_1 _10765_ (.A(net520),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__mux4_1 _10766_ (.A0(\dpath.RF.R[16][27] ),
    .A1(\dpath.RF.R[17][27] ),
    .A2(\dpath.RF.R[18][27] ),
    .A3(\dpath.RF.R[19][27] ),
    .S0(net575),
    .S1(net556),
    .X(_04957_));
 sky130_fd_sc_hd__nor2_1 _10767_ (.A(net536),
    .B(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__mux4_1 _10768_ (.A0(\dpath.RF.R[20][27] ),
    .A1(\dpath.RF.R[21][27] ),
    .A2(\dpath.RF.R[22][27] ),
    .A3(\dpath.RF.R[23][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04959_));
 sky130_fd_sc_hd__nor2_1 _10769_ (.A(net515),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__mux4_1 _10770_ (.A0(\dpath.RF.R[28][27] ),
    .A1(\dpath.RF.R[29][27] ),
    .A2(\dpath.RF.R[30][27] ),
    .A3(\dpath.RF.R[31][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04961_));
 sky130_fd_sc_hd__nor2_1 _10771_ (.A(net515),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__mux4_1 _10772_ (.A0(\dpath.RF.R[24][27] ),
    .A1(\dpath.RF.R[25][27] ),
    .A2(\dpath.RF.R[26][27] ),
    .A3(\dpath.RF.R[27][27] ),
    .S0(net573),
    .S1(net554),
    .X(_04963_));
 sky130_fd_sc_hd__o21ai_1 _10773_ (.A1(net536),
    .A2(_04963_),
    .B1(net526),
    .Y(_04964_));
 sky130_fd_sc_hd__o32a_1 _10774_ (.A1(net526),
    .A2(_04958_),
    .A3(_04960_),
    .B1(_04962_),
    .B2(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__a221o_1 _10775_ (.A1(_04951_),
    .A2(_04956_),
    .B1(_04965_),
    .B2(net520),
    .C1(net483),
    .X(_04966_));
 sky130_fd_sc_hd__nor2_1 _10776_ (.A(net371),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__mux2_2 _10777_ (.A0(net3667),
    .A1(net20),
    .S(net479),
    .X(_04968_));
 sky130_fd_sc_hd__a221o_1 _10778_ (.A1(net663),
    .A2(net369),
    .B1(net367),
    .B2(_04968_),
    .C1(_04967_),
    .X(_04969_));
 sky130_fd_sc_hd__a22oi_1 _10779_ (.A1(net648),
    .A2(\dpath.alu.adder.in1[26] ),
    .B1(\dpath.alu.adder.in1[27] ),
    .B2(net652),
    .Y(_04970_));
 sky130_fd_sc_hd__and3_1 _10780_ (.A(net652),
    .B(net648),
    .C(\dpath.alu.adder.in1[27] ),
    .X(_04971_));
 sky130_fd_sc_hd__and2_1 _10781_ (.A(\dpath.alu.adder.in1[26] ),
    .B(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__or2_1 _10782_ (.A(_04970_),
    .B(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__a22o_1 _10783_ (.A1(net640),
    .A2(net720),
    .B1(\dpath.alu.adder.in1[25] ),
    .B2(net644),
    .X(_04974_));
 sky130_fd_sc_hd__and3_1 _10784_ (.A(net644),
    .B(net640),
    .C(\dpath.alu.adder.in1[25] ),
    .X(_04975_));
 sky130_fd_sc_hd__a21bo_1 _10785_ (.A1(net720),
    .A2(_04975_),
    .B1_N(_04974_),
    .X(_04976_));
 sky130_fd_sc_hd__nand2_1 _10786_ (.A(net634),
    .B(net721),
    .Y(_04977_));
 sky130_fd_sc_hd__xnor2_1 _10787_ (.A(_04976_),
    .B(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__or2_1 _10788_ (.A(_04798_),
    .B(_04800_),
    .X(_04979_));
 sky130_fd_sc_hd__and2b_1 _10789_ (.A_N(_04978_),
    .B(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__xor2_1 _10790_ (.A(_04978_),
    .B(_04979_),
    .X(_04981_));
 sky130_fd_sc_hd__nor2_1 _10791_ (.A(_04973_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__xor2_1 _10792_ (.A(_04973_),
    .B(_04981_),
    .X(_04983_));
 sky130_fd_sc_hd__and2b_1 _10793_ (.A_N(_04805_),
    .B(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__xnor2_1 _10794_ (.A(_04805_),
    .B(_04983_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_1 _10795_ (.A(_04817_),
    .B(_04819_),
    .Y(_04986_));
 sky130_fd_sc_hd__a22o_1 _10796_ (.A1(net614),
    .A2(net728),
    .B1(net726),
    .B2(net618),
    .X(_04987_));
 sky130_fd_sc_hd__and4_1 _10797_ (.A(net618),
    .B(net614),
    .C(net728),
    .D(net726),
    .X(_04988_));
 sky130_fd_sc_hd__nand4_1 _10798_ (.A(net618),
    .B(net614),
    .C(net728),
    .D(net726),
    .Y(_04989_));
 sky130_fd_sc_hd__and2_1 _10799_ (.A(net610),
    .B(net730),
    .X(_04990_));
 sky130_fd_sc_hd__a21oi_1 _10800_ (.A1(_04987_),
    .A2(_04989_),
    .B1(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__and3_1 _10801_ (.A(_04987_),
    .B(_04989_),
    .C(_04990_),
    .X(_04992_));
 sky130_fd_sc_hd__nor2_1 _10802_ (.A(_04991_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__a22o_1 _10803_ (.A1(net626),
    .A2(net723),
    .B1(net722),
    .B2(net630),
    .X(_04994_));
 sky130_fd_sc_hd__nand4_2 _10804_ (.A(net630),
    .B(net626),
    .C(net723),
    .D(net722),
    .Y(_04995_));
 sky130_fd_sc_hd__inv_2 _10805_ (.A(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__a22oi_2 _10806_ (.A1(net622),
    .A2(net725),
    .B1(_04994_),
    .B2(_04995_),
    .Y(_04997_));
 sky130_fd_sc_hd__and4_2 _10807_ (.A(net622),
    .B(net725),
    .C(_04994_),
    .D(_04995_),
    .X(_04998_));
 sky130_fd_sc_hd__a211o_1 _10808_ (.A1(_04813_),
    .A2(_04815_),
    .B1(_04997_),
    .C1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__o211ai_2 _10809_ (.A1(_04997_),
    .A2(_04998_),
    .B1(_04813_),
    .C1(_04815_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand3_2 _10810_ (.A(_04993_),
    .B(_04999_),
    .C(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__a21o_1 _10811_ (.A1(_04999_),
    .A2(_05000_),
    .B1(_04993_),
    .X(_05002_));
 sky130_fd_sc_hd__nand3_4 _10812_ (.A(_04803_),
    .B(_05001_),
    .C(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__a21o_1 _10813_ (.A1(_05001_),
    .A2(_05002_),
    .B1(_04803_),
    .X(_05004_));
 sky130_fd_sc_hd__nand3_4 _10814_ (.A(_04986_),
    .B(_05003_),
    .C(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__a21o_1 _10815_ (.A1(_05003_),
    .A2(_05004_),
    .B1(_04986_),
    .X(_05006_));
 sky130_fd_sc_hd__and3_1 _10816_ (.A(_04985_),
    .B(_05005_),
    .C(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__nand3_1 _10817_ (.A(_04985_),
    .B(_05005_),
    .C(_05006_),
    .Y(_05008_));
 sky130_fd_sc_hd__a21o_1 _10818_ (.A1(_05005_),
    .A2(_05006_),
    .B1(_04985_),
    .X(_05009_));
 sky130_fd_sc_hd__nand3_2 _10819_ (.A(_04825_),
    .B(_05008_),
    .C(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__a21o_1 _10820_ (.A1(_05008_),
    .A2(_05009_),
    .B1(_04825_),
    .X(_05011_));
 sky130_fd_sc_hd__a22o_1 _10821_ (.A1(net753),
    .A2(net589),
    .B1(net587),
    .B2(net756),
    .X(_05012_));
 sky130_fd_sc_hd__and3_1 _10822_ (.A(net756),
    .B(net753),
    .C(net589),
    .X(_05013_));
 sky130_fd_sc_hd__a21bo_1 _10823_ (.A1(net587),
    .A2(_05013_),
    .B1_N(_05012_),
    .X(_05014_));
 sky130_fd_sc_hd__nand2_1 _10824_ (.A(net759),
    .B(net585),
    .Y(_05015_));
 sky130_fd_sc_hd__xor2_2 _10825_ (.A(_05014_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__and4_1 _10826_ (.A(net743),
    .B(net739),
    .C(net599),
    .D(net595),
    .X(_05017_));
 sky130_fd_sc_hd__nand4_1 _10827_ (.A(\dpath.alu.adder.in1[12] ),
    .B(net739),
    .C(net598),
    .D(net596),
    .Y(_05018_));
 sky130_fd_sc_hd__a22o_1 _10828_ (.A1(\dpath.alu.adder.in1[13] ),
    .A2(net598),
    .B1(net596),
    .B2(\dpath.alu.adder.in1[12] ),
    .X(_05019_));
 sky130_fd_sc_hd__and4_1 _10829_ (.A(net747),
    .B(net592),
    .C(_05018_),
    .D(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__nand4_1 _10830_ (.A(\dpath.alu.adder.in1[11] ),
    .B(net593),
    .C(_05018_),
    .D(_05019_),
    .Y(_05021_));
 sky130_fd_sc_hd__a22o_1 _10831_ (.A1(net747),
    .A2(net593),
    .B1(_05018_),
    .B2(_05019_),
    .X(_05022_));
 sky130_fd_sc_hd__o211a_1 _10832_ (.A1(_04834_),
    .A2(_04837_),
    .B1(_05021_),
    .C1(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__a211o_1 _10833_ (.A1(_05021_),
    .A2(_05022_),
    .B1(_04834_),
    .C1(_04837_),
    .X(_05024_));
 sky130_fd_sc_hd__nand2b_1 _10834_ (.A_N(_05023_),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__xnor2_2 _10835_ (.A(_05016_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _10836_ (.A(_04846_),
    .B(_04848_),
    .Y(_05027_));
 sky130_fd_sc_hd__nand4_2 _10837_ (.A(net607),
    .B(net605),
    .C(net735),
    .D(net733),
    .Y(_05028_));
 sky130_fd_sc_hd__inv_2 _10838_ (.A(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__a22o_1 _10839_ (.A1(net605),
    .A2(net735),
    .B1(net733),
    .B2(net607),
    .X(_05030_));
 sky130_fd_sc_hd__and4_1 _10840_ (.A(net602),
    .B(net738),
    .C(_05028_),
    .D(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__a22oi_2 _10841_ (.A1(net602),
    .A2(net738),
    .B1(_05028_),
    .B2(_05030_),
    .Y(_05032_));
 sky130_fd_sc_hd__a211o_1 _10842_ (.A1(_04809_),
    .A2(_04811_),
    .B1(_05031_),
    .C1(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__o211ai_2 _10843_ (.A1(_05031_),
    .A2(_05032_),
    .B1(_04809_),
    .C1(_04811_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand3_1 _10844_ (.A(_05027_),
    .B(_05033_),
    .C(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__a21o_1 _10845_ (.A1(_05033_),
    .A2(_05034_),
    .B1(_05027_),
    .X(_05036_));
 sky130_fd_sc_hd__a21bo_1 _10846_ (.A1(_04844_),
    .A2(_04851_),
    .B1_N(_04850_),
    .X(_05037_));
 sky130_fd_sc_hd__and3_1 _10847_ (.A(_05035_),
    .B(_05036_),
    .C(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__nand3_1 _10848_ (.A(_05035_),
    .B(_05036_),
    .C(_05037_),
    .Y(_05039_));
 sky130_fd_sc_hd__a21o_1 _10849_ (.A1(_05035_),
    .A2(_05036_),
    .B1(_05037_),
    .X(_05040_));
 sky130_fd_sc_hd__and3_2 _10850_ (.A(_05026_),
    .B(_05039_),
    .C(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__a21oi_2 _10851_ (.A1(_05039_),
    .A2(_05040_),
    .B1(_05026_),
    .Y(_05042_));
 sky130_fd_sc_hd__a211o_2 _10852_ (.A1(_04821_),
    .A2(_04823_),
    .B1(_05041_),
    .C1(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__o211ai_4 _10853_ (.A1(_05041_),
    .A2(_05042_),
    .B1(_04821_),
    .C1(_04823_),
    .Y(_05044_));
 sky130_fd_sc_hd__o211ai_4 _10854_ (.A1(_04855_),
    .A2(_04858_),
    .B1(_05043_),
    .C1(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__a211o_1 _10855_ (.A1(_05043_),
    .A2(_05044_),
    .B1(_04855_),
    .C1(_04858_),
    .X(_05046_));
 sky130_fd_sc_hd__nand4_2 _10856_ (.A(_05010_),
    .B(_05011_),
    .C(_05045_),
    .D(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__a22o_1 _10857_ (.A1(_05010_),
    .A2(_05011_),
    .B1(_05045_),
    .B2(_05046_),
    .X(_05048_));
 sky130_fd_sc_hd__o211a_1 _10858_ (.A1(_04827_),
    .A2(_04865_),
    .B1(_05047_),
    .C1(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__a211oi_1 _10859_ (.A1(_05047_),
    .A2(_05048_),
    .B1(_04827_),
    .C1(_04865_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand4_1 _10860_ (.A(net777),
    .B(net772),
    .C(net579),
    .D(\dpath.alu.adder.in0[24] ),
    .Y(_05051_));
 sky130_fd_sc_hd__a22o_1 _10861_ (.A1(net772),
    .A2(net579),
    .B1(\dpath.alu.adder.in0[24] ),
    .B2(net777),
    .X(_05052_));
 sky130_fd_sc_hd__and2_1 _10862_ (.A(net780),
    .B(\dpath.alu.adder.in0[25] ),
    .X(_05053_));
 sky130_fd_sc_hd__nand3_1 _10863_ (.A(_05051_),
    .B(_05052_),
    .C(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__a21o_1 _10864_ (.A1(_05051_),
    .A2(_05052_),
    .B1(_05053_),
    .X(_05055_));
 sky130_fd_sc_hd__a21bo_1 _10865_ (.A1(_04871_),
    .A2(_04872_),
    .B1_N(_04870_),
    .X(_05056_));
 sky130_fd_sc_hd__and3_1 _10866_ (.A(_05054_),
    .B(_05055_),
    .C(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__a21oi_1 _10867_ (.A1(_05054_),
    .A2(_05055_),
    .B1(_05056_),
    .Y(_05058_));
 sky130_fd_sc_hd__or2_1 _10868_ (.A(_05057_),
    .B(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__nand2_1 _10869_ (.A(net784),
    .B(\dpath.alu.adder.in0[26] ),
    .Y(_05060_));
 sky130_fd_sc_hd__xnor2_1 _10870_ (.A(_05059_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21ba_1 _10871_ (.A1(_04877_),
    .A2(_04879_),
    .B1_N(_04876_),
    .X(_05062_));
 sky130_fd_sc_hd__xor2_1 _10872_ (.A(_05061_),
    .B(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__and2_1 _10873_ (.A(net786),
    .B(\dpath.alu.adder.in0[27] ),
    .X(_05064_));
 sky130_fd_sc_hd__nor2_1 _10874_ (.A(_05063_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__and2_1 _10875_ (.A(_05063_),
    .B(_05064_),
    .X(_05066_));
 sky130_fd_sc_hd__or2_1 _10876_ (.A(_05065_),
    .B(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__a21o_1 _10877_ (.A1(_04833_),
    .A2(_04841_),
    .B1(_04840_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _10878_ (.A(_04890_),
    .B(_04892_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand4_1 _10879_ (.A(net764),
    .B(net760),
    .C(net583),
    .D(net581),
    .Y(_05070_));
 sky130_fd_sc_hd__a22o_1 _10880_ (.A1(net760),
    .A2(net583),
    .B1(net581),
    .B2(net764),
    .X(_05071_));
 sky130_fd_sc_hd__and4_1 _10881_ (.A(net768),
    .B(net580),
    .C(_05070_),
    .D(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__a22oi_2 _10882_ (.A1(net768),
    .A2(net580),
    .B1(_05070_),
    .B2(_05071_),
    .Y(_05073_));
 sky130_fd_sc_hd__a211o_2 _10883_ (.A1(_04829_),
    .A2(_04831_),
    .B1(_05072_),
    .C1(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__o211ai_2 _10884_ (.A1(_05072_),
    .A2(_05073_),
    .B1(_04829_),
    .C1(_04831_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand3_2 _10885_ (.A(_05069_),
    .B(_05074_),
    .C(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a21o_1 _10886_ (.A1(_05074_),
    .A2(_05075_),
    .B1(_05069_),
    .X(_05077_));
 sky130_fd_sc_hd__and3_2 _10887_ (.A(_05068_),
    .B(_05076_),
    .C(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a21oi_2 _10888_ (.A1(_05076_),
    .A2(_05077_),
    .B1(_05068_),
    .Y(_05079_));
 sky130_fd_sc_hd__a211oi_4 _10889_ (.A1(_04894_),
    .A2(_04896_),
    .B1(_05078_),
    .C1(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__o211a_1 _10890_ (.A1(_05078_),
    .A2(_05079_),
    .B1(_04894_),
    .C1(_04896_),
    .X(_05081_));
 sky130_fd_sc_hd__a211oi_2 _10891_ (.A1(_04899_),
    .A2(_04901_),
    .B1(_05080_),
    .C1(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__o211a_1 _10892_ (.A1(_05080_),
    .A2(_05081_),
    .B1(_04899_),
    .C1(_04901_),
    .X(_05083_));
 sky130_fd_sc_hd__or3_2 _10893_ (.A(_05067_),
    .B(_05082_),
    .C(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__o21ai_2 _10894_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_05067_),
    .Y(_05085_));
 sky130_fd_sc_hd__o211ai_2 _10895_ (.A1(_04861_),
    .A2(_04863_),
    .B1(_05084_),
    .C1(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__inv_2 _10896_ (.A(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__a211o_1 _10897_ (.A1(_05084_),
    .A2(_05085_),
    .B1(_04861_),
    .C1(_04863_),
    .X(_05088_));
 sky130_fd_sc_hd__o211a_1 _10898_ (.A1(_04903_),
    .A2(_04905_),
    .B1(_05086_),
    .C1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__a211oi_1 _10899_ (.A1(_05086_),
    .A2(_05088_),
    .B1(_04903_),
    .C1(_04905_),
    .Y(_05090_));
 sky130_fd_sc_hd__or4_2 _10900_ (.A(_05049_),
    .B(_05050_),
    .C(_05089_),
    .D(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__o22ai_2 _10901_ (.A1(_05049_),
    .A2(_05050_),
    .B1(_05089_),
    .B2(_05090_),
    .Y(_05092_));
 sky130_fd_sc_hd__o211a_1 _10902_ (.A1(_04867_),
    .A2(_04911_),
    .B1(_05091_),
    .C1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__a211oi_1 _10903_ (.A1(_05091_),
    .A2(_05092_),
    .B1(_04867_),
    .C1(_04911_),
    .Y(_05094_));
 sky130_fd_sc_hd__a211oi_2 _10904_ (.A1(_04907_),
    .A2(_04909_),
    .B1(_05093_),
    .C1(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__o211a_1 _10905_ (.A1(_05093_),
    .A2(_05094_),
    .B1(_04907_),
    .C1(_04909_),
    .X(_05096_));
 sky130_fd_sc_hd__a211oi_2 _10906_ (.A1(_04913_),
    .A2(_04915_),
    .B1(_05095_),
    .C1(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__o211a_1 _10907_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_04913_),
    .C1(_04915_),
    .X(_05098_));
 sky130_fd_sc_hd__a211oi_2 _10908_ (.A1(_04882_),
    .A2(_04885_),
    .B1(_05097_),
    .C1(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__o211a_1 _10909_ (.A1(_05097_),
    .A2(_05098_),
    .B1(_04882_),
    .C1(_04885_),
    .X(_05100_));
 sky130_fd_sc_hd__o211a_1 _10910_ (.A1(_05099_),
    .A2(_05100_),
    .B1(_04918_),
    .C1(_04920_),
    .X(_05101_));
 sky130_fd_sc_hd__a211o_1 _10911_ (.A1(_04918_),
    .A2(_04920_),
    .B1(_05099_),
    .C1(_05100_),
    .X(_05102_));
 sky130_fd_sc_hd__nand2b_1 _10912_ (.A_N(_05101_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__o21ai_1 _10913_ (.A1(_04926_),
    .A2(_04929_),
    .B1(_04924_),
    .Y(_05104_));
 sky130_fd_sc_hd__xnor2_1 _10914_ (.A(_05103_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(net3646),
    .A1(_05105_),
    .S(_02071_),
    .X(_05106_));
 sky130_fd_sc_hd__a21oi_1 _10916_ (.A1(_01915_),
    .A2(_04794_),
    .B1(_01875_),
    .Y(_05107_));
 sky130_fd_sc_hd__a31o_1 _10917_ (.A1(_01875_),
    .A2(_01915_),
    .A3(_04794_),
    .B1(net469),
    .X(_05108_));
 sky130_fd_sc_hd__a2bb2o_4 _10918_ (.A1_N(_05107_),
    .A2_N(_05108_),
    .B1(net469),
    .B2(_05106_),
    .X(_05109_));
 sky130_fd_sc_hd__a21oi_4 _10919_ (.A1(net391),
    .A2(_05109_),
    .B1(_04969_),
    .Y(_05110_));
 sky130_fd_sc_hd__nor2_1 _10920_ (.A(net374),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__xnor2_1 _10921_ (.A(net578),
    .B(net3339),
    .Y(_05112_));
 sky130_fd_sc_hd__o21a_1 _10922_ (.A1(_04937_),
    .A2(_04940_),
    .B1(_04936_),
    .X(_05113_));
 sky130_fd_sc_hd__xnor2_1 _10923_ (.A(_05112_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__nor2_1 _10924_ (.A(net366),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_1 _10925_ (.A(net247),
    .B(_04943_),
    .Y(_05116_));
 sky130_fd_sc_hd__o211a_1 _10926_ (.A1(net247),
    .A2(_04943_),
    .B1(_05116_),
    .C1(net362),
    .X(_05117_));
 sky130_fd_sc_hd__a2111o_1 _10927_ (.A1(net3252),
    .A2(net404),
    .B1(net451),
    .C1(_05115_),
    .D1(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__o221a_1 _10928_ (.A1(net247),
    .A2(net444),
    .B1(_05111_),
    .B2(net3253),
    .C1(net852),
    .X(_00663_));
 sky130_fd_sc_hd__mux4_1 _10929_ (.A0(\dpath.RF.R[0][28] ),
    .A1(\dpath.RF.R[1][28] ),
    .A2(\dpath.RF.R[2][28] ),
    .A3(\dpath.RF.R[3][28] ),
    .S0(net573),
    .S1(net554),
    .X(_05119_));
 sky130_fd_sc_hd__mux4_1 _10930_ (.A0(\dpath.RF.R[4][28] ),
    .A1(\dpath.RF.R[5][28] ),
    .A2(\dpath.RF.R[6][28] ),
    .A3(\dpath.RF.R[7][28] ),
    .S0(net573),
    .S1(net554),
    .X(_05120_));
 sky130_fd_sc_hd__o21a_1 _10931_ (.A1(net515),
    .A2(_05120_),
    .B1(net507),
    .X(_05121_));
 sky130_fd_sc_hd__o21ai_1 _10932_ (.A1(net536),
    .A2(_05119_),
    .B1(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__mux4_1 _10933_ (.A0(\dpath.RF.R[12][28] ),
    .A1(\dpath.RF.R[13][28] ),
    .A2(\dpath.RF.R[14][28] ),
    .A3(\dpath.RF.R[15][28] ),
    .S0(net574),
    .S1(net555),
    .X(_05123_));
 sky130_fd_sc_hd__mux4_1 _10934_ (.A0(\dpath.RF.R[8][28] ),
    .A1(\dpath.RF.R[9][28] ),
    .A2(\dpath.RF.R[10][28] ),
    .A3(\dpath.RF.R[11][28] ),
    .S0(net574),
    .S1(net555),
    .X(_05124_));
 sky130_fd_sc_hd__or2_1 _10935_ (.A(net536),
    .B(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__o211a_1 _10936_ (.A1(net515),
    .A2(_05123_),
    .B1(_05125_),
    .C1(net526),
    .X(_05126_));
 sky130_fd_sc_hd__nor2_1 _10937_ (.A(net520),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__mux4_1 _10938_ (.A0(\dpath.RF.R[16][28] ),
    .A1(\dpath.RF.R[17][28] ),
    .A2(\dpath.RF.R[18][28] ),
    .A3(\dpath.RF.R[19][28] ),
    .S0(net574),
    .S1(net555),
    .X(_05128_));
 sky130_fd_sc_hd__nor2_1 _10939_ (.A(net536),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__mux4_1 _10940_ (.A0(\dpath.RF.R[20][28] ),
    .A1(\dpath.RF.R[21][28] ),
    .A2(\dpath.RF.R[22][28] ),
    .A3(\dpath.RF.R[23][28] ),
    .S0(net574),
    .S1(net555),
    .X(_05130_));
 sky130_fd_sc_hd__nor2_1 _10941_ (.A(net515),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__mux4_1 _10942_ (.A0(\dpath.RF.R[28][28] ),
    .A1(\dpath.RF.R[29][28] ),
    .A2(\dpath.RF.R[30][28] ),
    .A3(\dpath.RF.R[31][28] ),
    .S0(net574),
    .S1(net555),
    .X(_05132_));
 sky130_fd_sc_hd__nor2_1 _10943_ (.A(net515),
    .B(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__mux4_1 _10944_ (.A0(\dpath.RF.R[24][28] ),
    .A1(\dpath.RF.R[25][28] ),
    .A2(\dpath.RF.R[26][28] ),
    .A3(\dpath.RF.R[27][28] ),
    .S0(net574),
    .S1(net555),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_1 _10945_ (.A1(net536),
    .A2(_05134_),
    .B1(net526),
    .Y(_05135_));
 sky130_fd_sc_hd__o32a_1 _10946_ (.A1(net526),
    .A2(_05129_),
    .A3(_05131_),
    .B1(_05133_),
    .B2(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__a221o_1 _10947_ (.A1(_05122_),
    .A2(_05127_),
    .B1(_05136_),
    .B2(net520),
    .C1(net483),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_1 _10948_ (.A(net371),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__mux2_2 _10949_ (.A0(net3676),
    .A1(net21),
    .S(net479),
    .X(_05139_));
 sky130_fd_sc_hd__a221o_1 _10950_ (.A1(net660),
    .A2(net370),
    .B1(net367),
    .B2(_05139_),
    .C1(_05138_),
    .X(_05140_));
 sky130_fd_sc_hd__or2_1 _10951_ (.A(_01875_),
    .B(_01916_),
    .X(_05141_));
 sky130_fd_sc_hd__or2_1 _10952_ (.A(_04792_),
    .B(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__a311o_1 _10953_ (.A1(_01918_),
    .A2(_01921_),
    .A3(_04272_),
    .B1(_05142_),
    .C1(_01917_),
    .X(_05143_));
 sky130_fd_sc_hd__o221a_1 _10954_ (.A1(_01873_),
    .A2(_01915_),
    .B1(_04791_),
    .B2(_05141_),
    .C1(_01874_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_1 _10955_ (.A(_05143_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__nor2_1 _10956_ (.A(_01938_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__a21o_1 _10957_ (.A1(_01938_),
    .A2(_05145_),
    .B1(net469),
    .X(_05147_));
 sky130_fd_sc_hd__or2_1 _10958_ (.A(_04926_),
    .B(_05103_),
    .X(_05148_));
 sky130_fd_sc_hd__a211o_1 _10959_ (.A1(_04458_),
    .A2(_04461_),
    .B1(_04928_),
    .C1(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__o221a_2 _10960_ (.A1(_04924_),
    .A2(_05101_),
    .B1(_05148_),
    .B2(_04927_),
    .C1(_05102_),
    .X(_05150_));
 sky130_fd_sc_hd__a22o_1 _10961_ (.A1(net648),
    .A2(\dpath.alu.adder.in1[27] ),
    .B1(\dpath.alu.adder.in1[28] ),
    .B2(net652),
    .X(_05151_));
 sky130_fd_sc_hd__a21bo_1 _10962_ (.A1(\dpath.alu.adder.in1[28] ),
    .A2(_04971_),
    .B1_N(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__nand2_1 _10963_ (.A(net644),
    .B(\dpath.alu.adder.in1[26] ),
    .Y(_05153_));
 sky130_fd_sc_hd__xor2_1 _10964_ (.A(_05152_),
    .B(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__a32o_1 _10965_ (.A1(net634),
    .A2(net721),
    .A3(_04974_),
    .B1(_04975_),
    .B2(net720),
    .X(_05155_));
 sky130_fd_sc_hd__a22o_1 _10966_ (.A1(net634),
    .A2(net720),
    .B1(\dpath.alu.adder.in1[25] ),
    .B2(net640),
    .X(_05156_));
 sky130_fd_sc_hd__nand4_2 _10967_ (.A(net640),
    .B(net634),
    .C(net720),
    .D(\dpath.alu.adder.in1[25] ),
    .Y(_05157_));
 sky130_fd_sc_hd__a22o_1 _10968_ (.A1(net630),
    .A2(net721),
    .B1(_05156_),
    .B2(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__nand4_2 _10969_ (.A(net630),
    .B(net721),
    .C(_05156_),
    .D(_05157_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand3_1 _10970_ (.A(_04972_),
    .B(_05158_),
    .C(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__a21o_1 _10971_ (.A1(_05158_),
    .A2(_05159_),
    .B1(_04972_),
    .X(_05161_));
 sky130_fd_sc_hd__nand3_1 _10972_ (.A(_05155_),
    .B(_05160_),
    .C(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__a21o_1 _10973_ (.A1(_05160_),
    .A2(_05161_),
    .B1(_05155_),
    .X(_05163_));
 sky130_fd_sc_hd__and3_1 _10974_ (.A(_05154_),
    .B(_05162_),
    .C(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__a21oi_1 _10975_ (.A1(_05162_),
    .A2(_05163_),
    .B1(_05154_),
    .Y(_05165_));
 sky130_fd_sc_hd__or3b_4 _10976_ (.A(_05164_),
    .B(_05165_),
    .C_N(_04982_),
    .X(_05166_));
 sky130_fd_sc_hd__o21bai_2 _10977_ (.A1(_05164_),
    .A2(_05165_),
    .B1_N(_04982_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_1 _10978_ (.A(_04999_),
    .B(_05001_),
    .Y(_05168_));
 sky130_fd_sc_hd__a22o_1 _10979_ (.A1(net610),
    .A2(net728),
    .B1(net726),
    .B2(net614),
    .X(_05169_));
 sky130_fd_sc_hd__and3_1 _10980_ (.A(net614),
    .B(net610),
    .C(net726),
    .X(_05170_));
 sky130_fd_sc_hd__a21bo_1 _10981_ (.A1(net728),
    .A2(_05170_),
    .B1_N(_05169_),
    .X(_05171_));
 sky130_fd_sc_hd__nand2_1 _10982_ (.A(net607),
    .B(net730),
    .Y(_05172_));
 sky130_fd_sc_hd__xor2_1 _10983_ (.A(_05171_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__a22o_1 _10984_ (.A1(net622),
    .A2(net723),
    .B1(net722),
    .B2(net626),
    .X(_05174_));
 sky130_fd_sc_hd__nand4_4 _10985_ (.A(net626),
    .B(net622),
    .C(net723),
    .D(net722),
    .Y(_05175_));
 sky130_fd_sc_hd__a22o_1 _10986_ (.A1(net618),
    .A2(net725),
    .B1(_05174_),
    .B2(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__nand4_4 _10987_ (.A(net618),
    .B(net725),
    .C(_05174_),
    .D(_05175_),
    .Y(_05177_));
 sky130_fd_sc_hd__o211ai_4 _10988_ (.A1(_04996_),
    .A2(_04998_),
    .B1(_05176_),
    .C1(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a211o_1 _10989_ (.A1(_05176_),
    .A2(_05177_),
    .B1(_04996_),
    .C1(_04998_),
    .X(_05179_));
 sky130_fd_sc_hd__nand3_2 _10990_ (.A(_05173_),
    .B(_05178_),
    .C(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__a21o_1 _10991_ (.A1(_05178_),
    .A2(_05179_),
    .B1(_05173_),
    .X(_05181_));
 sky130_fd_sc_hd__nand3_2 _10992_ (.A(_04980_),
    .B(_05180_),
    .C(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__a21o_1 _10993_ (.A1(_05180_),
    .A2(_05181_),
    .B1(_04980_),
    .X(_05183_));
 sky130_fd_sc_hd__nand3_2 _10994_ (.A(_05168_),
    .B(_05182_),
    .C(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__a21o_1 _10995_ (.A1(_05182_),
    .A2(_05183_),
    .B1(_05168_),
    .X(_05185_));
 sky130_fd_sc_hd__nand4_4 _10996_ (.A(_05166_),
    .B(_05167_),
    .C(_05184_),
    .D(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__a22o_1 _10997_ (.A1(_05166_),
    .A2(_05167_),
    .B1(_05184_),
    .B2(_05185_),
    .X(_05187_));
 sky130_fd_sc_hd__o211ai_4 _10998_ (.A1(_04984_),
    .A2(_05007_),
    .B1(_05186_),
    .C1(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__a211o_1 _10999_ (.A1(_05186_),
    .A2(_05187_),
    .B1(_04984_),
    .C1(_05007_),
    .X(_05189_));
 sky130_fd_sc_hd__a22o_1 _11000_ (.A1(net753),
    .A2(net587),
    .B1(net585),
    .B2(net756),
    .X(_05190_));
 sky130_fd_sc_hd__and3_1 _11001_ (.A(net756),
    .B(net753),
    .C(net587),
    .X(_05191_));
 sky130_fd_sc_hd__a21bo_1 _11002_ (.A1(net585),
    .A2(_05191_),
    .B1_N(_05190_),
    .X(_05192_));
 sky130_fd_sc_hd__nand2_1 _11003_ (.A(net759),
    .B(net583),
    .Y(_05193_));
 sky130_fd_sc_hd__xor2_2 _11004_ (.A(_05192_),
    .B(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__a22o_1 _11005_ (.A1(net739),
    .A2(net595),
    .B1(net592),
    .B2(net743),
    .X(_05195_));
 sky130_fd_sc_hd__and4_1 _11006_ (.A(net743),
    .B(net739),
    .C(net595),
    .D(net592),
    .X(_05196_));
 sky130_fd_sc_hd__nand4_1 _11007_ (.A(net743),
    .B(net739),
    .C(net595),
    .D(net592),
    .Y(_05197_));
 sky130_fd_sc_hd__a22o_1 _11008_ (.A1(net747),
    .A2(net589),
    .B1(_05195_),
    .B2(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__and4_1 _11009_ (.A(net747),
    .B(net589),
    .C(_05195_),
    .D(_05197_),
    .X(_05199_));
 sky130_fd_sc_hd__nand4_1 _11010_ (.A(net747),
    .B(net589),
    .C(_05195_),
    .D(_05197_),
    .Y(_05200_));
 sky130_fd_sc_hd__o211a_1 _11011_ (.A1(_05017_),
    .A2(_05020_),
    .B1(_05198_),
    .C1(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__a211o_1 _11012_ (.A1(_05198_),
    .A2(_05200_),
    .B1(_05017_),
    .C1(_05020_),
    .X(_05202_));
 sky130_fd_sc_hd__nand2b_1 _11013_ (.A_N(_05201_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__xnor2_2 _11014_ (.A(_05194_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__or2_1 _11015_ (.A(_05029_),
    .B(_05031_),
    .X(_05205_));
 sky130_fd_sc_hd__a22o_1 _11016_ (.A1(net602),
    .A2(net735),
    .B1(net733),
    .B2(net605),
    .X(_05206_));
 sky130_fd_sc_hd__nand4_2 _11017_ (.A(net605),
    .B(net602),
    .C(net735),
    .D(net733),
    .Y(_05207_));
 sky130_fd_sc_hd__nand3b_2 _11018_ (.A_N(_01895_),
    .B(_05206_),
    .C(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__a21bo_1 _11019_ (.A1(_05206_),
    .A2(_05207_),
    .B1_N(_01895_),
    .X(_05209_));
 sky130_fd_sc_hd__o211ai_2 _11020_ (.A1(_04988_),
    .A2(_04992_),
    .B1(_05208_),
    .C1(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__a211o_1 _11021_ (.A1(_05208_),
    .A2(_05209_),
    .B1(_04988_),
    .C1(_04992_),
    .X(_05211_));
 sky130_fd_sc_hd__nand3_1 _11022_ (.A(_05205_),
    .B(_05210_),
    .C(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__a21o_1 _11023_ (.A1(_05210_),
    .A2(_05211_),
    .B1(_05205_),
    .X(_05213_));
 sky130_fd_sc_hd__a21bo_1 _11024_ (.A1(_05027_),
    .A2(_05034_),
    .B1_N(_05033_),
    .X(_05214_));
 sky130_fd_sc_hd__and3_1 _11025_ (.A(_05212_),
    .B(_05213_),
    .C(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__a21oi_1 _11026_ (.A1(_05212_),
    .A2(_05213_),
    .B1(_05214_),
    .Y(_05216_));
 sky130_fd_sc_hd__nor3b_2 _11027_ (.A(_05215_),
    .B(_05216_),
    .C_N(_05204_),
    .Y(_05217_));
 sky130_fd_sc_hd__o21ba_1 _11028_ (.A1(_05215_),
    .A2(_05216_),
    .B1_N(_05204_),
    .X(_05218_));
 sky130_fd_sc_hd__a211o_2 _11029_ (.A1(_05003_),
    .A2(_05005_),
    .B1(_05217_),
    .C1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__o211ai_4 _11030_ (.A1(_05217_),
    .A2(_05218_),
    .B1(_05003_),
    .C1(_05005_),
    .Y(_05220_));
 sky130_fd_sc_hd__o211ai_4 _11031_ (.A1(_05038_),
    .A2(_05041_),
    .B1(_05219_),
    .C1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__a211o_1 _11032_ (.A1(_05219_),
    .A2(_05220_),
    .B1(_05038_),
    .C1(_05041_),
    .X(_05222_));
 sky130_fd_sc_hd__nand4_2 _11033_ (.A(_05188_),
    .B(_05189_),
    .C(_05221_),
    .D(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a22o_1 _11034_ (.A1(_05188_),
    .A2(_05189_),
    .B1(_05221_),
    .B2(_05222_),
    .X(_05224_));
 sky130_fd_sc_hd__nand2_1 _11035_ (.A(_05223_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__a21o_1 _11036_ (.A1(_05010_),
    .A2(_05047_),
    .B1(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__nand3_1 _11037_ (.A(_05010_),
    .B(_05047_),
    .C(_05225_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand2b_2 _11038_ (.A_N(_05082_),
    .B(_05084_),
    .Y(_05228_));
 sky130_fd_sc_hd__inv_2 _11039_ (.A(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__nand4_2 _11040_ (.A(net777),
    .B(net775),
    .C(\dpath.alu.adder.in0[24] ),
    .D(\dpath.alu.adder.in0[25] ),
    .Y(_05230_));
 sky130_fd_sc_hd__a22o_1 _11041_ (.A1(net775),
    .A2(\dpath.alu.adder.in0[24] ),
    .B1(\dpath.alu.adder.in0[25] ),
    .B2(net777),
    .X(_05231_));
 sky130_fd_sc_hd__nand4_2 _11042_ (.A(net780),
    .B(\dpath.alu.adder.in0[26] ),
    .C(_05230_),
    .D(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__a22o_1 _11043_ (.A1(net780),
    .A2(\dpath.alu.adder.in0[26] ),
    .B1(_05230_),
    .B2(_05231_),
    .X(_05233_));
 sky130_fd_sc_hd__a21bo_1 _11044_ (.A1(_05052_),
    .A2(_05053_),
    .B1_N(_05051_),
    .X(_05234_));
 sky130_fd_sc_hd__and3_1 _11045_ (.A(_05232_),
    .B(_05233_),
    .C(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__a21oi_1 _11046_ (.A1(_05232_),
    .A2(_05233_),
    .B1(_05234_),
    .Y(_05236_));
 sky130_fd_sc_hd__or2_1 _11047_ (.A(_05235_),
    .B(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__nand2_1 _11048_ (.A(net784),
    .B(\dpath.alu.adder.in0[27] ),
    .Y(_05238_));
 sky130_fd_sc_hd__xnor2_1 _11049_ (.A(_05237_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__o21ba_1 _11050_ (.A1(_05058_),
    .A2(_05060_),
    .B1_N(_05057_),
    .X(_05240_));
 sky130_fd_sc_hd__or2_1 _11051_ (.A(_05239_),
    .B(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__xor2_1 _11052_ (.A(_05239_),
    .B(_05240_),
    .X(_05242_));
 sky130_fd_sc_hd__nand2_1 _11053_ (.A(net787),
    .B(\dpath.alu.adder.in0[28] ),
    .Y(_05243_));
 sky130_fd_sc_hd__nand3_1 _11054_ (.A(net787),
    .B(\dpath.alu.adder.in0[28] ),
    .C(_05242_),
    .Y(_05244_));
 sky130_fd_sc_hd__xor2_1 _11055_ (.A(_05242_),
    .B(_05243_),
    .X(_05245_));
 sky130_fd_sc_hd__a21o_1 _11056_ (.A1(_05016_),
    .A2(_05024_),
    .B1(_05023_),
    .X(_05246_));
 sky130_fd_sc_hd__a41o_1 _11057_ (.A1(net764),
    .A2(net760),
    .A3(net583),
    .A4(net581),
    .B1(_05072_),
    .X(_05247_));
 sky130_fd_sc_hd__a32o_1 _11058_ (.A1(net759),
    .A2(net585),
    .A3(_05012_),
    .B1(_05013_),
    .B2(net587),
    .X(_05248_));
 sky130_fd_sc_hd__a22o_1 _11059_ (.A1(net760),
    .A2(net581),
    .B1(net580),
    .B2(net764),
    .X(_05249_));
 sky130_fd_sc_hd__nand4_2 _11060_ (.A(net764),
    .B(net760),
    .C(net581),
    .D(net580),
    .Y(_05250_));
 sky130_fd_sc_hd__a22o_1 _11061_ (.A1(net768),
    .A2(net579),
    .B1(_05249_),
    .B2(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__nand4_2 _11062_ (.A(net768),
    .B(net579),
    .C(_05249_),
    .D(_05250_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand3_1 _11063_ (.A(_05248_),
    .B(_05251_),
    .C(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__a21o_1 _11064_ (.A1(_05251_),
    .A2(_05252_),
    .B1(_05248_),
    .X(_05254_));
 sky130_fd_sc_hd__nand3_1 _11065_ (.A(_05247_),
    .B(_05253_),
    .C(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__a21o_1 _11066_ (.A1(_05253_),
    .A2(_05254_),
    .B1(_05247_),
    .X(_05256_));
 sky130_fd_sc_hd__and3_2 _11067_ (.A(_05246_),
    .B(_05255_),
    .C(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__a21oi_2 _11068_ (.A1(_05255_),
    .A2(_05256_),
    .B1(_05246_),
    .Y(_05258_));
 sky130_fd_sc_hd__a211oi_2 _11069_ (.A1(_05074_),
    .A2(_05076_),
    .B1(_05257_),
    .C1(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__a211o_1 _11070_ (.A1(_05074_),
    .A2(_05076_),
    .B1(_05257_),
    .C1(_05258_),
    .X(_05260_));
 sky130_fd_sc_hd__o211ai_2 _11071_ (.A1(_05257_),
    .A2(_05258_),
    .B1(_05074_),
    .C1(_05076_),
    .Y(_05261_));
 sky130_fd_sc_hd__o211a_1 _11072_ (.A1(_05078_),
    .A2(_05080_),
    .B1(_05260_),
    .C1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__inv_2 _11073_ (.A(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__a211oi_2 _11074_ (.A1(_05260_),
    .A2(_05261_),
    .B1(_05078_),
    .C1(_05080_),
    .Y(_05264_));
 sky130_fd_sc_hd__nor3_1 _11075_ (.A(_05245_),
    .B(_05262_),
    .C(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__or3_1 _11076_ (.A(_05245_),
    .B(_05262_),
    .C(_05264_),
    .X(_05266_));
 sky130_fd_sc_hd__o21a_1 _11077_ (.A1(_05262_),
    .A2(_05264_),
    .B1(_05245_),
    .X(_05267_));
 sky130_fd_sc_hd__a211oi_1 _11078_ (.A1(_05043_),
    .A2(_05045_),
    .B1(_05265_),
    .C1(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__o211a_1 _11079_ (.A1(_05265_),
    .A2(_05267_),
    .B1(_05043_),
    .C1(_05045_),
    .X(_05269_));
 sky130_fd_sc_hd__or2_1 _11080_ (.A(_05268_),
    .B(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__xnor2_2 _11081_ (.A(_05228_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand3_2 _11082_ (.A(_05226_),
    .B(_05227_),
    .C(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__a21o_1 _11083_ (.A1(_05226_),
    .A2(_05227_),
    .B1(_05271_),
    .X(_05273_));
 sky130_fd_sc_hd__nand2_1 _11084_ (.A(_05272_),
    .B(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2b_1 _11085_ (.A_N(_05049_),
    .B(_05091_),
    .Y(_05275_));
 sky130_fd_sc_hd__and3_1 _11086_ (.A(_05272_),
    .B(_05273_),
    .C(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__xnor2_1 _11087_ (.A(_05274_),
    .B(_05275_),
    .Y(_05277_));
 sky130_fd_sc_hd__o21a_1 _11088_ (.A1(_05087_),
    .A2(_05089_),
    .B1(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__or3_1 _11089_ (.A(_05087_),
    .B(_05089_),
    .C(_05277_),
    .X(_05279_));
 sky130_fd_sc_hd__and2b_1 _11090_ (.A_N(_05278_),
    .B(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__nor2_1 _11091_ (.A(_05093_),
    .B(_05095_),
    .Y(_05281_));
 sky130_fd_sc_hd__and2b_1 _11092_ (.A_N(_05281_),
    .B(_05280_),
    .X(_05282_));
 sky130_fd_sc_hd__xnor2_1 _11093_ (.A(_05280_),
    .B(_05281_),
    .Y(_05283_));
 sky130_fd_sc_hd__o21bai_2 _11094_ (.A1(_05061_),
    .A2(_05062_),
    .B1_N(_05066_),
    .Y(_05284_));
 sky130_fd_sc_hd__and2_1 _11095_ (.A(_05283_),
    .B(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__xnor2_1 _11096_ (.A(_05283_),
    .B(_05284_),
    .Y(_05286_));
 sky130_fd_sc_hd__o21ba_2 _11097_ (.A1(_05097_),
    .A2(_05099_),
    .B1_N(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__or3b_1 _11098_ (.A(_05097_),
    .B(_05099_),
    .C_N(_05286_),
    .X(_05288_));
 sky130_fd_sc_hd__nand2b_1 _11099_ (.A_N(_05287_),
    .B(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__a21oi_4 _11100_ (.A1(_05149_),
    .A2(_05150_),
    .B1(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__a311o_1 _11101_ (.A1(_05149_),
    .A2(_05150_),
    .A3(_05289_),
    .B1(_05290_),
    .C1(_02240_),
    .X(_05291_));
 sky130_fd_sc_hd__o221ai_4 _11102_ (.A1(_01787_),
    .A2(net484),
    .B1(_05146_),
    .B2(_05147_),
    .C1(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__a21o_2 _11103_ (.A1(net391),
    .A2(_05292_),
    .B1(_05140_),
    .X(_05293_));
 sky130_fd_sc_hd__and2_1 _11104_ (.A(_02027_),
    .B(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__or2_1 _11105_ (.A(net578),
    .B(net3401),
    .X(_05295_));
 sky130_fd_sc_hd__nand2_1 _11106_ (.A(net578),
    .B(net3401),
    .Y(_05296_));
 sky130_fd_sc_hd__nand2_1 _11107_ (.A(_05295_),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__or4_1 _11108_ (.A(_04597_),
    .B(_04937_),
    .C(_04938_),
    .D(_05112_),
    .X(_05298_));
 sky130_fd_sc_hd__o21a_1 _11109_ (.A1(net3339),
    .A2(net3509),
    .B1(net578),
    .X(_05299_));
 sky130_fd_sc_hd__nor2_1 _11110_ (.A(_04939_),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _11111_ (.A(_05298_),
    .B(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__xor2_1 _11112_ (.A(_05297_),
    .B(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__and3_1 _11113_ (.A(net3471),
    .B(net3441),
    .C(_04943_),
    .X(_05303_));
 sky130_fd_sc_hd__a21oi_1 _11114_ (.A1(net3441),
    .A2(_04943_),
    .B1(net3471),
    .Y(_05304_));
 sky130_fd_sc_hd__a21oi_1 _11115_ (.A1(\dpath.btarg_DX.q[28] ),
    .A2(net404),
    .B1(net451),
    .Y(_05305_));
 sky130_fd_sc_hd__o31a_1 _11116_ (.A1(_01958_),
    .A2(_05303_),
    .A3(_05304_),
    .B1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__o21ai_1 _11117_ (.A1(net366),
    .A2(_05302_),
    .B1(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__o221a_1 _11118_ (.A1(net3471),
    .A2(net444),
    .B1(_05294_),
    .B2(_05307_),
    .C1(net858),
    .X(_00664_));
 sky130_fd_sc_hd__mux4_1 _11119_ (.A0(\dpath.RF.R[0][29] ),
    .A1(\dpath.RF.R[1][29] ),
    .A2(\dpath.RF.R[2][29] ),
    .A3(\dpath.RF.R[3][29] ),
    .S0(net575),
    .S1(net556),
    .X(_05308_));
 sky130_fd_sc_hd__mux4_1 _11120_ (.A0(\dpath.RF.R[4][29] ),
    .A1(\dpath.RF.R[5][29] ),
    .A2(\dpath.RF.R[6][29] ),
    .A3(\dpath.RF.R[7][29] ),
    .S0(net574),
    .S1(net555),
    .X(_05309_));
 sky130_fd_sc_hd__o21a_1 _11121_ (.A1(net516),
    .A2(_05309_),
    .B1(net507),
    .X(_05310_));
 sky130_fd_sc_hd__o21ai_1 _11122_ (.A1(net537),
    .A2(_05308_),
    .B1(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__mux4_1 _11123_ (.A0(\dpath.RF.R[12][29] ),
    .A1(\dpath.RF.R[13][29] ),
    .A2(\dpath.RF.R[14][29] ),
    .A3(\dpath.RF.R[15][29] ),
    .S0(net575),
    .S1(net556),
    .X(_05312_));
 sky130_fd_sc_hd__mux4_1 _11124_ (.A0(\dpath.RF.R[8][29] ),
    .A1(\dpath.RF.R[9][29] ),
    .A2(\dpath.RF.R[10][29] ),
    .A3(\dpath.RF.R[11][29] ),
    .S0(net575),
    .S1(net556),
    .X(_05313_));
 sky130_fd_sc_hd__or2_1 _11125_ (.A(net537),
    .B(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__o211a_1 _11126_ (.A1(net516),
    .A2(_05312_),
    .B1(_05314_),
    .C1(net526),
    .X(_05315_));
 sky130_fd_sc_hd__nor2_1 _11127_ (.A(net520),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__mux4_1 _11128_ (.A0(\dpath.RF.R[16][29] ),
    .A1(\dpath.RF.R[17][29] ),
    .A2(\dpath.RF.R[18][29] ),
    .A3(\dpath.RF.R[19][29] ),
    .S0(net574),
    .S1(net555),
    .X(_05317_));
 sky130_fd_sc_hd__nor2_1 _11129_ (.A(net536),
    .B(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__mux4_1 _11130_ (.A0(\dpath.RF.R[20][29] ),
    .A1(\dpath.RF.R[21][29] ),
    .A2(\dpath.RF.R[22][29] ),
    .A3(\dpath.RF.R[23][29] ),
    .S0(net574),
    .S1(net555),
    .X(_05319_));
 sky130_fd_sc_hd__nor2_1 _11131_ (.A(net515),
    .B(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__mux4_1 _11132_ (.A0(\dpath.RF.R[28][29] ),
    .A1(\dpath.RF.R[29][29] ),
    .A2(\dpath.RF.R[30][29] ),
    .A3(\dpath.RF.R[31][29] ),
    .S0(net574),
    .S1(net555),
    .X(_05321_));
 sky130_fd_sc_hd__nor2_1 _11133_ (.A(net515),
    .B(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__mux4_1 _11134_ (.A0(\dpath.RF.R[24][29] ),
    .A1(\dpath.RF.R[25][29] ),
    .A2(\dpath.RF.R[26][29] ),
    .A3(\dpath.RF.R[27][29] ),
    .S0(net574),
    .S1(net555),
    .X(_05323_));
 sky130_fd_sc_hd__o21ai_1 _11135_ (.A1(net536),
    .A2(_05323_),
    .B1(net526),
    .Y(_05324_));
 sky130_fd_sc_hd__o32a_1 _11136_ (.A1(net526),
    .A2(_05318_),
    .A3(_05320_),
    .B1(_05322_),
    .B2(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__a221o_1 _11137_ (.A1(_05311_),
    .A2(_05316_),
    .B1(_05325_),
    .B2(net520),
    .C1(net483),
    .X(_05326_));
 sky130_fd_sc_hd__nor2_1 _11138_ (.A(net371),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__mux2_2 _11139_ (.A0(net3663),
    .A1(net22),
    .S(net480),
    .X(_05328_));
 sky130_fd_sc_hd__a221o_1 _11140_ (.A1(net659),
    .A2(net369),
    .B1(net367),
    .B2(_05328_),
    .C1(_05327_),
    .X(_05329_));
 sky130_fd_sc_hd__nand2_1 _11141_ (.A(net652),
    .B(\dpath.alu.adder.in1[29] ),
    .Y(_05330_));
 sky130_fd_sc_hd__a22o_1 _11142_ (.A1(net644),
    .A2(\dpath.alu.adder.in1[27] ),
    .B1(\dpath.alu.adder.in1[28] ),
    .B2(net648),
    .X(_05331_));
 sky130_fd_sc_hd__nand4_1 _11143_ (.A(net648),
    .B(net644),
    .C(\dpath.alu.adder.in1[27] ),
    .D(\dpath.alu.adder.in1[28] ),
    .Y(_05332_));
 sky130_fd_sc_hd__and2_1 _11144_ (.A(net640),
    .B(\dpath.alu.adder.in1[26] ),
    .X(_05333_));
 sky130_fd_sc_hd__a21oi_1 _11145_ (.A1(_05331_),
    .A2(_05332_),
    .B1(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__and3_1 _11146_ (.A(_05331_),
    .B(_05332_),
    .C(_05333_),
    .X(_05335_));
 sky130_fd_sc_hd__nor2_1 _11147_ (.A(_05334_),
    .B(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__nor3_1 _11148_ (.A(_05330_),
    .B(_05334_),
    .C(_05335_),
    .Y(_05337_));
 sky130_fd_sc_hd__xnor2_1 _11149_ (.A(_05330_),
    .B(_05336_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _11150_ (.A(_05157_),
    .B(_05159_),
    .Y(_05339_));
 sky130_fd_sc_hd__a32o_1 _11151_ (.A1(net644),
    .A2(\dpath.alu.adder.in1[26] ),
    .A3(_05151_),
    .B1(_04971_),
    .B2(\dpath.alu.adder.in1[28] ),
    .X(_05340_));
 sky130_fd_sc_hd__a22o_1 _11152_ (.A1(net630),
    .A2(net720),
    .B1(\dpath.alu.adder.in1[25] ),
    .B2(net634),
    .X(_05341_));
 sky130_fd_sc_hd__nand4_2 _11153_ (.A(net634),
    .B(net630),
    .C(net720),
    .D(\dpath.alu.adder.in1[25] ),
    .Y(_05342_));
 sky130_fd_sc_hd__a22o_1 _11154_ (.A1(net626),
    .A2(net721),
    .B1(_05341_),
    .B2(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__nand4_2 _11155_ (.A(net626),
    .B(net721),
    .C(_05341_),
    .D(_05342_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand3_1 _11156_ (.A(_05340_),
    .B(_05343_),
    .C(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__a21o_1 _11157_ (.A1(_05343_),
    .A2(_05344_),
    .B1(_05340_),
    .X(_05346_));
 sky130_fd_sc_hd__nand3_1 _11158_ (.A(_05339_),
    .B(_05345_),
    .C(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__a21o_1 _11159_ (.A1(_05345_),
    .A2(_05346_),
    .B1(_05339_),
    .X(_05348_));
 sky130_fd_sc_hd__and3_1 _11160_ (.A(_05338_),
    .B(_05347_),
    .C(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__a21oi_1 _11161_ (.A1(_05347_),
    .A2(_05348_),
    .B1(_05338_),
    .Y(_05350_));
 sky130_fd_sc_hd__nor3b_2 _11162_ (.A(_05349_),
    .B(_05350_),
    .C_N(_05164_),
    .Y(_05351_));
 sky130_fd_sc_hd__o21ba_1 _11163_ (.A1(_05349_),
    .A2(_05350_),
    .B1_N(_05164_),
    .X(_05352_));
 sky130_fd_sc_hd__a21bo_1 _11164_ (.A1(_05155_),
    .A2(_05161_),
    .B1_N(_05160_),
    .X(_05353_));
 sky130_fd_sc_hd__a22o_1 _11165_ (.A1(net607),
    .A2(net728),
    .B1(net726),
    .B2(net610),
    .X(_05354_));
 sky130_fd_sc_hd__and3_1 _11166_ (.A(net610),
    .B(net607),
    .C(net726),
    .X(_05355_));
 sky130_fd_sc_hd__a21bo_1 _11167_ (.A1(net728),
    .A2(_05355_),
    .B1_N(_05354_),
    .X(_05356_));
 sky130_fd_sc_hd__nand2_1 _11168_ (.A(net604),
    .B(net730),
    .Y(_05357_));
 sky130_fd_sc_hd__xor2_1 _11169_ (.A(_05356_),
    .B(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__a22o_1 _11170_ (.A1(net618),
    .A2(net723),
    .B1(net722),
    .B2(net622),
    .X(_05359_));
 sky130_fd_sc_hd__nand4_1 _11171_ (.A(net622),
    .B(net618),
    .C(net723),
    .D(net722),
    .Y(_05360_));
 sky130_fd_sc_hd__and2_1 _11172_ (.A(net614),
    .B(net725),
    .X(_05361_));
 sky130_fd_sc_hd__a21oi_1 _11173_ (.A1(_05359_),
    .A2(_05360_),
    .B1(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__and3_1 _11174_ (.A(_05359_),
    .B(_05360_),
    .C(_05361_),
    .X(_05363_));
 sky130_fd_sc_hd__a211o_1 _11175_ (.A1(_05175_),
    .A2(_05177_),
    .B1(_05362_),
    .C1(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__o211ai_2 _11176_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05175_),
    .C1(_05177_),
    .Y(_05365_));
 sky130_fd_sc_hd__nand3_2 _11177_ (.A(_05358_),
    .B(_05364_),
    .C(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__a21o_1 _11178_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05358_),
    .X(_05367_));
 sky130_fd_sc_hd__and3_1 _11179_ (.A(_05353_),
    .B(_05366_),
    .C(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__a21oi_1 _11180_ (.A1(_05366_),
    .A2(_05367_),
    .B1(_05353_),
    .Y(_05369_));
 sky130_fd_sc_hd__a211oi_2 _11181_ (.A1(_05178_),
    .A2(_05180_),
    .B1(_05368_),
    .C1(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__o211a_1 _11182_ (.A1(_05368_),
    .A2(_05369_),
    .B1(_05178_),
    .C1(_05180_),
    .X(_05371_));
 sky130_fd_sc_hd__nor4_2 _11183_ (.A(_05351_),
    .B(_05352_),
    .C(_05370_),
    .D(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__o22a_1 _11184_ (.A1(_05351_),
    .A2(_05352_),
    .B1(_05370_),
    .B2(_05371_),
    .X(_05373_));
 sky130_fd_sc_hd__a211o_1 _11185_ (.A1(_05166_),
    .A2(_05186_),
    .B1(_05372_),
    .C1(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__inv_2 _11186_ (.A(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__o211ai_2 _11187_ (.A1(_05372_),
    .A2(_05373_),
    .B1(_05166_),
    .C1(_05186_),
    .Y(_05376_));
 sky130_fd_sc_hd__a22o_1 _11188_ (.A1(net753),
    .A2(net585),
    .B1(net583),
    .B2(net756),
    .X(_05377_));
 sky130_fd_sc_hd__and3_1 _11189_ (.A(net756),
    .B(net753),
    .C(net585),
    .X(_05378_));
 sky130_fd_sc_hd__a21bo_1 _11190_ (.A1(net583),
    .A2(_05378_),
    .B1_N(_05377_),
    .X(_05379_));
 sky130_fd_sc_hd__nand2_1 _11191_ (.A(net759),
    .B(net581),
    .Y(_05380_));
 sky130_fd_sc_hd__xor2_1 _11192_ (.A(_05379_),
    .B(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__a22o_1 _11193_ (.A1(net739),
    .A2(net592),
    .B1(net589),
    .B2(net743),
    .X(_05382_));
 sky130_fd_sc_hd__nand4_2 _11194_ (.A(net743),
    .B(net739),
    .C(net592),
    .D(net589),
    .Y(_05383_));
 sky130_fd_sc_hd__a22o_1 _11195_ (.A1(net747),
    .A2(net587),
    .B1(_05382_),
    .B2(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__nand4_2 _11196_ (.A(net747),
    .B(net587),
    .C(_05382_),
    .D(_05383_),
    .Y(_05385_));
 sky130_fd_sc_hd__o211a_1 _11197_ (.A1(_05196_),
    .A2(_05199_),
    .B1(_05384_),
    .C1(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__a211o_1 _11198_ (.A1(_05384_),
    .A2(_05385_),
    .B1(_05196_),
    .C1(_05199_),
    .X(_05387_));
 sky130_fd_sc_hd__nand2b_1 _11199_ (.A_N(_05386_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__xnor2_1 _11200_ (.A(_05381_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(_05207_),
    .B(_05208_),
    .Y(_05390_));
 sky130_fd_sc_hd__a32o_1 _11202_ (.A1(net609),
    .A2(net730),
    .A3(_05169_),
    .B1(_05170_),
    .B2(net728),
    .X(_05391_));
 sky130_fd_sc_hd__a22o_1 _11203_ (.A1(net599),
    .A2(net735),
    .B1(net733),
    .B2(net602),
    .X(_05392_));
 sky130_fd_sc_hd__nand4_1 _11204_ (.A(net602),
    .B(net599),
    .C(net735),
    .D(net733),
    .Y(_05393_));
 sky130_fd_sc_hd__a22o_1 _11205_ (.A1(net738),
    .A2(net595),
    .B1(_05392_),
    .B2(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__nand4_1 _11206_ (.A(net738),
    .B(net595),
    .C(_05392_),
    .D(_05393_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand3_1 _11207_ (.A(_05391_),
    .B(_05394_),
    .C(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__a21o_1 _11208_ (.A1(_05394_),
    .A2(_05395_),
    .B1(_05391_),
    .X(_05397_));
 sky130_fd_sc_hd__nand3_1 _11209_ (.A(_05390_),
    .B(_05396_),
    .C(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__a21o_1 _11210_ (.A1(_05396_),
    .A2(_05397_),
    .B1(_05390_),
    .X(_05399_));
 sky130_fd_sc_hd__a21bo_1 _11211_ (.A1(_05205_),
    .A2(_05211_),
    .B1_N(_05210_),
    .X(_05400_));
 sky130_fd_sc_hd__and3_1 _11212_ (.A(_05398_),
    .B(_05399_),
    .C(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__a21oi_1 _11213_ (.A1(_05398_),
    .A2(_05399_),
    .B1(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__nor3b_2 _11214_ (.A(_05401_),
    .B(_05402_),
    .C_N(_05389_),
    .Y(_05403_));
 sky130_fd_sc_hd__o21ba_1 _11215_ (.A1(_05401_),
    .A2(_05402_),
    .B1_N(_05389_),
    .X(_05404_));
 sky130_fd_sc_hd__a211o_1 _11216_ (.A1(_05182_),
    .A2(_05184_),
    .B1(_05403_),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__o211ai_2 _11217_ (.A1(_05403_),
    .A2(_05404_),
    .B1(_05182_),
    .C1(_05184_),
    .Y(_05406_));
 sky130_fd_sc_hd__o211ai_2 _11218_ (.A1(_05215_),
    .A2(_05217_),
    .B1(_05405_),
    .C1(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__a211o_1 _11219_ (.A1(_05405_),
    .A2(_05406_),
    .B1(_05215_),
    .C1(_05217_),
    .X(_05408_));
 sky130_fd_sc_hd__and4_1 _11220_ (.A(_05374_),
    .B(_05376_),
    .C(_05407_),
    .D(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__a22oi_2 _11221_ (.A1(_05374_),
    .A2(_05376_),
    .B1(_05407_),
    .B2(_05408_),
    .Y(_05410_));
 sky130_fd_sc_hd__a211oi_2 _11222_ (.A1(_05188_),
    .A2(_05223_),
    .B1(_05409_),
    .C1(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__o211a_1 _11223_ (.A1(_05409_),
    .A2(_05410_),
    .B1(_05188_),
    .C1(_05223_),
    .X(_05412_));
 sky130_fd_sc_hd__a22oi_1 _11224_ (.A1(net775),
    .A2(\dpath.alu.adder.in0[25] ),
    .B1(\dpath.alu.adder.in0[26] ),
    .B2(net777),
    .Y(_05413_));
 sky130_fd_sc_hd__and4_1 _11225_ (.A(net777),
    .B(net775),
    .C(\dpath.alu.adder.in0[25] ),
    .D(\dpath.alu.adder.in0[26] ),
    .X(_05414_));
 sky130_fd_sc_hd__o2bb2a_1 _11226_ (.A1_N(net780),
    .A2_N(\dpath.alu.adder.in0[27] ),
    .B1(_05413_),
    .B2(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__and4bb_1 _11227_ (.A_N(_05413_),
    .B_N(_05414_),
    .C(net782),
    .D(\dpath.alu.adder.in0[27] ),
    .X(_05416_));
 sky130_fd_sc_hd__or2_1 _11228_ (.A(_05415_),
    .B(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__nand2_1 _11229_ (.A(_05230_),
    .B(_05232_),
    .Y(_05418_));
 sky130_fd_sc_hd__and2b_1 _11230_ (.A_N(_05417_),
    .B(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__xnor2_1 _11231_ (.A(_05417_),
    .B(_05418_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand2_1 _11232_ (.A(net784),
    .B(\dpath.alu.adder.in0[28] ),
    .Y(_05421_));
 sky130_fd_sc_hd__and3_1 _11233_ (.A(net784),
    .B(\dpath.alu.adder.in0[28] ),
    .C(_05420_),
    .X(_05422_));
 sky130_fd_sc_hd__xor2_1 _11234_ (.A(_05420_),
    .B(_05421_),
    .X(_05423_));
 sky130_fd_sc_hd__o21ba_1 _11235_ (.A1(_05236_),
    .A2(_05238_),
    .B1_N(_05235_),
    .X(_05424_));
 sky130_fd_sc_hd__xor2_1 _11236_ (.A(_05423_),
    .B(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(net787),
    .B(\dpath.alu.adder.in0[29] ),
    .Y(_05426_));
 sky130_fd_sc_hd__and3_1 _11238_ (.A(net787),
    .B(\dpath.alu.adder.in0[29] ),
    .C(_05425_),
    .X(_05427_));
 sky130_fd_sc_hd__xor2_1 _11239_ (.A(_05425_),
    .B(_05426_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _11240_ (.A(_05253_),
    .B(_05255_),
    .Y(_05429_));
 sky130_fd_sc_hd__a21o_1 _11241_ (.A1(_05194_),
    .A2(_05202_),
    .B1(_05201_),
    .X(_05430_));
 sky130_fd_sc_hd__nand2_1 _11242_ (.A(_05250_),
    .B(_05252_),
    .Y(_05431_));
 sky130_fd_sc_hd__a32o_1 _11243_ (.A1(net759),
    .A2(net583),
    .A3(_05190_),
    .B1(_05191_),
    .B2(net585),
    .X(_05432_));
 sky130_fd_sc_hd__a22o_1 _11244_ (.A1(net760),
    .A2(net580),
    .B1(net579),
    .B2(net764),
    .X(_05433_));
 sky130_fd_sc_hd__nand4_2 _11245_ (.A(net764),
    .B(net760),
    .C(net580),
    .D(net579),
    .Y(_05434_));
 sky130_fd_sc_hd__a22o_1 _11246_ (.A1(net768),
    .A2(\dpath.alu.adder.in0[24] ),
    .B1(_05433_),
    .B2(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__nand4_2 _11247_ (.A(net768),
    .B(\dpath.alu.adder.in0[24] ),
    .C(_05433_),
    .D(_05434_),
    .Y(_05436_));
 sky130_fd_sc_hd__nand3_2 _11248_ (.A(_05432_),
    .B(_05435_),
    .C(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21o_1 _11249_ (.A1(_05435_),
    .A2(_05436_),
    .B1(_05432_),
    .X(_05438_));
 sky130_fd_sc_hd__nand3_2 _11250_ (.A(_05431_),
    .B(_05437_),
    .C(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__a21o_1 _11251_ (.A1(_05437_),
    .A2(_05438_),
    .B1(_05431_),
    .X(_05440_));
 sky130_fd_sc_hd__nand3_2 _11252_ (.A(_05430_),
    .B(_05439_),
    .C(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__a21o_1 _11253_ (.A1(_05439_),
    .A2(_05440_),
    .B1(_05430_),
    .X(_05442_));
 sky130_fd_sc_hd__nand3_2 _11254_ (.A(_05429_),
    .B(_05441_),
    .C(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__a21o_1 _11255_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05429_),
    .X(_05444_));
 sky130_fd_sc_hd__o211a_1 _11256_ (.A1(_05257_),
    .A2(_05259_),
    .B1(_05443_),
    .C1(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__a211oi_2 _11257_ (.A1(_05443_),
    .A2(_05444_),
    .B1(_05257_),
    .C1(_05259_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor3_1 _11258_ (.A(_05428_),
    .B(_05445_),
    .C(_05446_),
    .Y(_05447_));
 sky130_fd_sc_hd__o21a_1 _11259_ (.A1(_05445_),
    .A2(_05446_),
    .B1(_05428_),
    .X(_05448_));
 sky130_fd_sc_hd__a211oi_2 _11260_ (.A1(_05219_),
    .A2(_05221_),
    .B1(_05447_),
    .C1(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__o211a_1 _11261_ (.A1(_05447_),
    .A2(_05448_),
    .B1(_05219_),
    .C1(_05221_),
    .X(_05450_));
 sky130_fd_sc_hd__a211oi_2 _11262_ (.A1(_05263_),
    .A2(_05266_),
    .B1(_05449_),
    .C1(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__o211a_1 _11263_ (.A1(_05449_),
    .A2(_05450_),
    .B1(_05263_),
    .C1(_05266_),
    .X(_05452_));
 sky130_fd_sc_hd__nor4_1 _11264_ (.A(_05411_),
    .B(_05412_),
    .C(_05451_),
    .D(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__o22a_1 _11265_ (.A1(_05411_),
    .A2(_05412_),
    .B1(_05451_),
    .B2(_05452_),
    .X(_05454_));
 sky130_fd_sc_hd__a211oi_2 _11266_ (.A1(_05226_),
    .A2(_05272_),
    .B1(net356),
    .C1(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__o211a_1 _11267_ (.A1(net356),
    .A2(_05454_),
    .B1(_05226_),
    .C1(_05272_),
    .X(_05456_));
 sky130_fd_sc_hd__o21ba_1 _11268_ (.A1(_05229_),
    .A2(_05270_),
    .B1_N(_05268_),
    .X(_05457_));
 sky130_fd_sc_hd__nor3_1 _11269_ (.A(_05455_),
    .B(_05456_),
    .C(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21a_1 _11270_ (.A1(_05455_),
    .A2(_05456_),
    .B1(_05457_),
    .X(_05459_));
 sky130_fd_sc_hd__nor2_1 _11271_ (.A(_05458_),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__o21a_1 _11272_ (.A1(_05276_),
    .A2(_05278_),
    .B1(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__nor3_1 _11273_ (.A(_05276_),
    .B(_05278_),
    .C(_05460_),
    .Y(_05462_));
 sky130_fd_sc_hd__a211oi_1 _11274_ (.A1(_05241_),
    .A2(_05244_),
    .B1(_05461_),
    .C1(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__o211a_1 _11275_ (.A1(_05461_),
    .A2(_05462_),
    .B1(_05241_),
    .C1(_05244_),
    .X(_05464_));
 sky130_fd_sc_hd__nor2_1 _11276_ (.A(_05463_),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__o21a_1 _11277_ (.A1(_05282_),
    .A2(_05285_),
    .B1(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__nor3_1 _11278_ (.A(_05282_),
    .B(_05285_),
    .C(_05465_),
    .Y(_05467_));
 sky130_fd_sc_hd__inv_2 _11279_ (.A(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__nor2_1 _11280_ (.A(_05466_),
    .B(_05467_),
    .Y(_05469_));
 sky130_fd_sc_hd__nor2_1 _11281_ (.A(_05287_),
    .B(_05290_),
    .Y(_05470_));
 sky130_fd_sc_hd__xnor2_1 _11282_ (.A(_05469_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__mux2_1 _11283_ (.A0(net3674),
    .A1(_05471_),
    .S(_02071_),
    .X(_05472_));
 sky130_fd_sc_hd__a21bo_1 _11284_ (.A1(_05143_),
    .A2(_05144_),
    .B1_N(_01936_),
    .X(_05473_));
 sky130_fd_sc_hd__nand2_1 _11285_ (.A(_01937_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__xor2_1 _11286_ (.A(_01860_),
    .B(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_2 _11287_ (.A0(_05472_),
    .A1(_05475_),
    .S(_02101_),
    .X(_05476_));
 sky130_fd_sc_hd__a21oi_4 _11288_ (.A1(net391),
    .A2(net3675),
    .B1(_05329_),
    .Y(_05477_));
 sky130_fd_sc_hd__nor2_1 _11289_ (.A(net374),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__nor2_1 _11290_ (.A(net578),
    .B(net3439),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _11291_ (.A(net578),
    .B(net3439),
    .Y(_05480_));
 sky130_fd_sc_hd__and2b_1 _11292_ (.A_N(_05479_),
    .B(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__a21bo_1 _11293_ (.A1(_05295_),
    .A2(_05301_),
    .B1_N(_05296_),
    .X(_05482_));
 sky130_fd_sc_hd__xnor2_1 _11294_ (.A(_05481_),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__and2_1 _11295_ (.A(net3447),
    .B(_05303_),
    .X(_05484_));
 sky130_fd_sc_hd__o21ai_1 _11296_ (.A1(net3447),
    .A2(_05303_),
    .B1(net362),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2_1 _11297_ (.A(net3491),
    .B(_01952_),
    .Y(_05486_));
 sky130_fd_sc_hd__o211a_1 _11298_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05486_),
    .C1(net444),
    .X(_05487_));
 sky130_fd_sc_hd__o21ai_1 _11299_ (.A1(net366),
    .A2(_05483_),
    .B1(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__o221a_1 _11300_ (.A1(net3447),
    .A2(net444),
    .B1(_05478_),
    .B2(_05488_),
    .C1(net858),
    .X(_00665_));
 sky130_fd_sc_hd__mux4_1 _11301_ (.A0(\dpath.RF.R[0][30] ),
    .A1(\dpath.RF.R[1][30] ),
    .A2(\dpath.RF.R[2][30] ),
    .A3(\dpath.RF.R[3][30] ),
    .S0(net571),
    .S1(net552),
    .X(_05489_));
 sky130_fd_sc_hd__mux4_1 _11302_ (.A0(\dpath.RF.R[4][30] ),
    .A1(\dpath.RF.R[5][30] ),
    .A2(\dpath.RF.R[6][30] ),
    .A3(\dpath.RF.R[7][30] ),
    .S0(net571),
    .S1(net552),
    .X(_05490_));
 sky130_fd_sc_hd__o21a_1 _11303_ (.A1(net516),
    .A2(_05490_),
    .B1(net507),
    .X(_05491_));
 sky130_fd_sc_hd__o21ai_1 _11304_ (.A1(net537),
    .A2(_05489_),
    .B1(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__mux4_1 _11305_ (.A0(\dpath.RF.R[12][30] ),
    .A1(\dpath.RF.R[13][30] ),
    .A2(\dpath.RF.R[14][30] ),
    .A3(\dpath.RF.R[15][30] ),
    .S0(net571),
    .S1(net552),
    .X(_05493_));
 sky130_fd_sc_hd__mux4_1 _11306_ (.A0(\dpath.RF.R[8][30] ),
    .A1(\dpath.RF.R[9][30] ),
    .A2(\dpath.RF.R[10][30] ),
    .A3(\dpath.RF.R[11][30] ),
    .S0(net571),
    .S1(net552),
    .X(_05494_));
 sky130_fd_sc_hd__or2_1 _11307_ (.A(net537),
    .B(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__o211a_1 _11308_ (.A1(net516),
    .A2(_05493_),
    .B1(_05495_),
    .C1(net527),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_1 _11309_ (.A(net520),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__mux4_1 _11310_ (.A0(\dpath.RF.R[16][30] ),
    .A1(\dpath.RF.R[17][30] ),
    .A2(\dpath.RF.R[18][30] ),
    .A3(\dpath.RF.R[19][30] ),
    .S0(net572),
    .S1(net553),
    .X(_05498_));
 sky130_fd_sc_hd__nor2_1 _11311_ (.A(net537),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__mux4_1 _11312_ (.A0(\dpath.RF.R[20][30] ),
    .A1(\dpath.RF.R[21][30] ),
    .A2(\dpath.RF.R[22][30] ),
    .A3(\dpath.RF.R[23][30] ),
    .S0(net572),
    .S1(net553),
    .X(_05500_));
 sky130_fd_sc_hd__nor2_1 _11313_ (.A(net516),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__mux4_1 _11314_ (.A0(\dpath.RF.R[28][30] ),
    .A1(\dpath.RF.R[29][30] ),
    .A2(\dpath.RF.R[30][30] ),
    .A3(\dpath.RF.R[31][30] ),
    .S0(net572),
    .S1(net553),
    .X(_05502_));
 sky130_fd_sc_hd__nor2_1 _11315_ (.A(net516),
    .B(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__mux4_1 _11316_ (.A0(\dpath.RF.R[24][30] ),
    .A1(\dpath.RF.R[25][30] ),
    .A2(\dpath.RF.R[26][30] ),
    .A3(\dpath.RF.R[27][30] ),
    .S0(net572),
    .S1(net553),
    .X(_05504_));
 sky130_fd_sc_hd__o21ai_1 _11317_ (.A1(net537),
    .A2(_05504_),
    .B1(net527),
    .Y(_05505_));
 sky130_fd_sc_hd__o32a_1 _11318_ (.A1(net527),
    .A2(_05499_),
    .A3(_05501_),
    .B1(_05503_),
    .B2(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__a221o_1 _11319_ (.A1(_05492_),
    .A2(_05497_),
    .B1(_05506_),
    .B2(net520),
    .C1(net483),
    .X(_05507_));
 sky130_fd_sc_hd__nor2_1 _11320_ (.A(net371),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__mux2_4 _11321_ (.A0(net3681),
    .A1(net24),
    .S(net480),
    .X(_05509_));
 sky130_fd_sc_hd__a221o_1 _11322_ (.A1(net656),
    .A2(_02115_),
    .B1(_02116_),
    .B2(_05509_),
    .C1(_05508_),
    .X(_05510_));
 sky130_fd_sc_hd__a21bo_1 _11323_ (.A1(_01937_),
    .A2(_05473_),
    .B1_N(_01858_),
    .X(_05511_));
 sky130_fd_sc_hd__a21o_1 _11324_ (.A1(_01859_),
    .A2(_05511_),
    .B1(_01884_),
    .X(_05512_));
 sky130_fd_sc_hd__a31oi_1 _11325_ (.A1(_01859_),
    .A2(_01884_),
    .A3(_05511_),
    .B1(net469),
    .Y(_05513_));
 sky130_fd_sc_hd__o31a_1 _11326_ (.A1(_05287_),
    .A2(_05290_),
    .A3(_05466_),
    .B1(_05468_),
    .X(_05514_));
 sky130_fd_sc_hd__o21ba_1 _11327_ (.A1(_05423_),
    .A2(_05424_),
    .B1_N(_05427_),
    .X(_05515_));
 sky130_fd_sc_hd__nor2_1 _11328_ (.A(_05449_),
    .B(_05451_),
    .Y(_05516_));
 sky130_fd_sc_hd__or2_1 _11329_ (.A(_05445_),
    .B(_05447_),
    .X(_05517_));
 sky130_fd_sc_hd__inv_2 _11330_ (.A(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__nand2_1 _11331_ (.A(_05405_),
    .B(_05407_),
    .Y(_05519_));
 sky130_fd_sc_hd__a22oi_1 _11332_ (.A1(net775),
    .A2(\dpath.alu.adder.in0[26] ),
    .B1(\dpath.alu.adder.in0[27] ),
    .B2(net777),
    .Y(_05520_));
 sky130_fd_sc_hd__and4_1 _11333_ (.A(net777),
    .B(net775),
    .C(\dpath.alu.adder.in0[26] ),
    .D(\dpath.alu.adder.in0[27] ),
    .X(_05521_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(_05520_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_1 _11335_ (.A(net782),
    .B(\dpath.alu.adder.in0[28] ),
    .Y(_05523_));
 sky130_fd_sc_hd__xor2_1 _11336_ (.A(_05522_),
    .B(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__or2_1 _11337_ (.A(_05414_),
    .B(_05416_),
    .X(_05525_));
 sky130_fd_sc_hd__and2b_1 _11338_ (.A_N(_05524_),
    .B(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__xor2_1 _11339_ (.A(_05524_),
    .B(_05525_),
    .X(_05527_));
 sky130_fd_sc_hd__nand2_1 _11340_ (.A(net784),
    .B(\dpath.alu.adder.in0[29] ),
    .Y(_05528_));
 sky130_fd_sc_hd__xor2_1 _11341_ (.A(_05527_),
    .B(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__o21a_1 _11342_ (.A1(_05419_),
    .A2(_05422_),
    .B1(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__nor3_1 _11343_ (.A(_05419_),
    .B(_05422_),
    .C(_05529_),
    .Y(_05531_));
 sky130_fd_sc_hd__nor2_1 _11344_ (.A(_05530_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _11345_ (.A(net787),
    .B(\dpath.alu.adder.in0[30] ),
    .Y(_05533_));
 sky130_fd_sc_hd__xor2_1 _11346_ (.A(_05532_),
    .B(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__a21o_1 _11347_ (.A1(_05381_),
    .A2(_05387_),
    .B1(_05386_),
    .X(_05535_));
 sky130_fd_sc_hd__nand2_1 _11348_ (.A(_05434_),
    .B(_05436_),
    .Y(_05536_));
 sky130_fd_sc_hd__a32o_1 _11349_ (.A1(net759),
    .A2(net581),
    .A3(_05377_),
    .B1(_05378_),
    .B2(net583),
    .X(_05537_));
 sky130_fd_sc_hd__a22o_1 _11350_ (.A1(net760),
    .A2(net579),
    .B1(\dpath.alu.adder.in0[24] ),
    .B2(net764),
    .X(_05538_));
 sky130_fd_sc_hd__nand4_1 _11351_ (.A(net764),
    .B(net760),
    .C(net579),
    .D(\dpath.alu.adder.in0[24] ),
    .Y(_05539_));
 sky130_fd_sc_hd__nand4_2 _11352_ (.A(net768),
    .B(\dpath.alu.adder.in0[25] ),
    .C(_05538_),
    .D(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__a22o_1 _11353_ (.A1(net768),
    .A2(\dpath.alu.adder.in0[25] ),
    .B1(_05538_),
    .B2(_05539_),
    .X(_05541_));
 sky130_fd_sc_hd__nand3_1 _11354_ (.A(_05537_),
    .B(_05540_),
    .C(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__a21o_1 _11355_ (.A1(_05540_),
    .A2(_05541_),
    .B1(_05537_),
    .X(_05543_));
 sky130_fd_sc_hd__nand3_1 _11356_ (.A(_05536_),
    .B(_05542_),
    .C(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__a21o_1 _11357_ (.A1(_05542_),
    .A2(_05543_),
    .B1(_05536_),
    .X(_05545_));
 sky130_fd_sc_hd__and3_1 _11358_ (.A(_05535_),
    .B(_05544_),
    .C(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__a21oi_1 _11359_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05535_),
    .Y(_05547_));
 sky130_fd_sc_hd__a211oi_2 _11360_ (.A1(_05437_),
    .A2(_05439_),
    .B1(_05546_),
    .C1(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__o211a_1 _11361_ (.A1(_05546_),
    .A2(_05547_),
    .B1(_05437_),
    .C1(_05439_),
    .X(_05549_));
 sky130_fd_sc_hd__a211oi_1 _11362_ (.A1(_05441_),
    .A2(_05443_),
    .B1(_05548_),
    .C1(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__o211a_1 _11363_ (.A1(_05548_),
    .A2(_05549_),
    .B1(_05441_),
    .C1(_05443_),
    .X(_05551_));
 sky130_fd_sc_hd__nor2_1 _11364_ (.A(_05550_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__xnor2_1 _11365_ (.A(_05534_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__and2_1 _11366_ (.A(_05519_),
    .B(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__xnor2_1 _11367_ (.A(_05519_),
    .B(_05553_),
    .Y(_05555_));
 sky130_fd_sc_hd__nor2_1 _11368_ (.A(_05518_),
    .B(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__xnor2_1 _11369_ (.A(_05518_),
    .B(_05555_),
    .Y(_05557_));
 sky130_fd_sc_hd__nor2_1 _11370_ (.A(_05401_),
    .B(_05403_),
    .Y(_05558_));
 sky130_fd_sc_hd__nor2_1 _11371_ (.A(_05368_),
    .B(_05370_),
    .Y(_05559_));
 sky130_fd_sc_hd__a22oi_1 _11372_ (.A1(net753),
    .A2(net583),
    .B1(net581),
    .B2(net756),
    .Y(_05560_));
 sky130_fd_sc_hd__and4_1 _11373_ (.A(net756),
    .B(net753),
    .C(net583),
    .D(net581),
    .X(_05561_));
 sky130_fd_sc_hd__nor2_1 _11374_ (.A(_05560_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _11375_ (.A(net759),
    .B(net580),
    .Y(_05563_));
 sky130_fd_sc_hd__xor2_1 _11376_ (.A(_05562_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__a22o_1 _11377_ (.A1(net739),
    .A2(net589),
    .B1(net587),
    .B2(net743),
    .X(_05565_));
 sky130_fd_sc_hd__nand4_1 _11378_ (.A(net743),
    .B(net739),
    .C(net589),
    .D(net587),
    .Y(_05566_));
 sky130_fd_sc_hd__nand2_1 _11379_ (.A(_05565_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand2_1 _11380_ (.A(net747),
    .B(net585),
    .Y(_05568_));
 sky130_fd_sc_hd__xor2_1 _11381_ (.A(_05567_),
    .B(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__nand2_1 _11382_ (.A(_05383_),
    .B(_05385_),
    .Y(_05570_));
 sky130_fd_sc_hd__xnor2_1 _11383_ (.A(_05569_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__nor2_1 _11384_ (.A(_05564_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__xor2_1 _11385_ (.A(_05564_),
    .B(_05571_),
    .X(_05573_));
 sky130_fd_sc_hd__nand2_1 _11386_ (.A(_05393_),
    .B(_05395_),
    .Y(_05574_));
 sky130_fd_sc_hd__a32o_1 _11387_ (.A1(net604),
    .A2(net730),
    .A3(_05354_),
    .B1(_05355_),
    .B2(net728),
    .X(_05575_));
 sky130_fd_sc_hd__a22o_1 _11388_ (.A1(net595),
    .A2(net735),
    .B1(net733),
    .B2(net599),
    .X(_05576_));
 sky130_fd_sc_hd__nand4_1 _11389_ (.A(net599),
    .B(net595),
    .C(net735),
    .D(net733),
    .Y(_05577_));
 sky130_fd_sc_hd__nand4_2 _11390_ (.A(net738),
    .B(net592),
    .C(_05576_),
    .D(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__a22o_1 _11391_ (.A1(net738),
    .A2(net592),
    .B1(_05576_),
    .B2(_05577_),
    .X(_05579_));
 sky130_fd_sc_hd__nand3_2 _11392_ (.A(_05575_),
    .B(_05578_),
    .C(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__a21o_1 _11393_ (.A1(_05578_),
    .A2(_05579_),
    .B1(_05575_),
    .X(_05581_));
 sky130_fd_sc_hd__nand3_2 _11394_ (.A(_05574_),
    .B(_05580_),
    .C(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__a21o_1 _11395_ (.A1(_05580_),
    .A2(_05581_),
    .B1(_05574_),
    .X(_05583_));
 sky130_fd_sc_hd__a21bo_1 _11396_ (.A1(_05390_),
    .A2(_05397_),
    .B1_N(_05396_),
    .X(_05584_));
 sky130_fd_sc_hd__nand3_1 _11397_ (.A(_05582_),
    .B(_05583_),
    .C(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__a21o_1 _11398_ (.A1(_05582_),
    .A2(_05583_),
    .B1(_05584_),
    .X(_05586_));
 sky130_fd_sc_hd__and3_1 _11399_ (.A(_05573_),
    .B(_05585_),
    .C(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__a21oi_1 _11400_ (.A1(_05585_),
    .A2(_05586_),
    .B1(_05573_),
    .Y(_05588_));
 sky130_fd_sc_hd__nor2_1 _11401_ (.A(_05587_),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__xnor2_1 _11402_ (.A(_05559_),
    .B(_05589_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand2b_1 _11403_ (.A_N(_05558_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__xnor2_1 _11404_ (.A(_05558_),
    .B(_05590_),
    .Y(_05592_));
 sky130_fd_sc_hd__a21bo_1 _11405_ (.A1(_05339_),
    .A2(_05346_),
    .B1_N(_05345_),
    .X(_05593_));
 sky130_fd_sc_hd__a22oi_1 _11406_ (.A1(net604),
    .A2(net728),
    .B1(net726),
    .B2(net609),
    .Y(_05594_));
 sky130_fd_sc_hd__and4_1 _11407_ (.A(net609),
    .B(net605),
    .C(net728),
    .D(net726),
    .X(_05595_));
 sky130_fd_sc_hd__nor2_1 _11408_ (.A(_05594_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(net602),
    .B(net730),
    .Y(_05597_));
 sky130_fd_sc_hd__xnor2_1 _11410_ (.A(_05596_),
    .B(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__a22o_1 _11411_ (.A1(net614),
    .A2(net723),
    .B1(net722),
    .B2(net618),
    .X(_05599_));
 sky130_fd_sc_hd__nand4_2 _11412_ (.A(net618),
    .B(net614),
    .C(net723),
    .D(net722),
    .Y(_05600_));
 sky130_fd_sc_hd__a22o_1 _11413_ (.A1(net610),
    .A2(net725),
    .B1(_05599_),
    .B2(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__nand4_2 _11414_ (.A(net610),
    .B(net725),
    .C(_05599_),
    .D(_05600_),
    .Y(_05602_));
 sky130_fd_sc_hd__a21bo_1 _11415_ (.A1(_05359_),
    .A2(_05361_),
    .B1_N(_05360_),
    .X(_05603_));
 sky130_fd_sc_hd__nand3_1 _11416_ (.A(_05601_),
    .B(_05602_),
    .C(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__a21o_1 _11417_ (.A1(_05601_),
    .A2(_05602_),
    .B1(_05603_),
    .X(_05605_));
 sky130_fd_sc_hd__nand3_1 _11418_ (.A(_05598_),
    .B(_05604_),
    .C(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__a21o_1 _11419_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05598_),
    .X(_05607_));
 sky130_fd_sc_hd__and3_1 _11420_ (.A(_05593_),
    .B(_05606_),
    .C(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__a21oi_1 _11421_ (.A1(_05606_),
    .A2(_05607_),
    .B1(_05593_),
    .Y(_05609_));
 sky130_fd_sc_hd__a211oi_2 _11422_ (.A1(_05364_),
    .A2(_05366_),
    .B1(_05608_),
    .C1(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__o211a_1 _11423_ (.A1(_05608_),
    .A2(_05609_),
    .B1(_05364_),
    .C1(_05366_),
    .X(_05611_));
 sky130_fd_sc_hd__a22o_1 _11424_ (.A1(net640),
    .A2(\dpath.alu.adder.in1[27] ),
    .B1(\dpath.alu.adder.in1[28] ),
    .B2(net644),
    .X(_05612_));
 sky130_fd_sc_hd__nand4_2 _11425_ (.A(net644),
    .B(net640),
    .C(\dpath.alu.adder.in1[27] ),
    .D(\dpath.alu.adder.in1[28] ),
    .Y(_05613_));
 sky130_fd_sc_hd__a22o_1 _11426_ (.A1(net634),
    .A2(\dpath.alu.adder.in1[26] ),
    .B1(_05612_),
    .B2(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__nand4_2 _11427_ (.A(net634),
    .B(\dpath.alu.adder.in1[26] ),
    .C(_05612_),
    .D(_05613_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_1 _11428_ (.A(net652),
    .B(\dpath.alu.adder.in1[30] ),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _11429_ (.A(net648),
    .B(\dpath.alu.adder.in1[29] ),
    .Y(_05617_));
 sky130_fd_sc_hd__xor2_1 _11430_ (.A(_05616_),
    .B(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__nand3_1 _11431_ (.A(_05614_),
    .B(_05615_),
    .C(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__a21o_1 _11432_ (.A1(_05614_),
    .A2(_05615_),
    .B1(_05618_),
    .X(_05620_));
 sky130_fd_sc_hd__a21oi_1 _11433_ (.A1(_05619_),
    .A2(_05620_),
    .B1(_05337_),
    .Y(_05621_));
 sky130_fd_sc_hd__and3_1 _11434_ (.A(_05337_),
    .B(_05619_),
    .C(_05620_),
    .X(_05622_));
 sky130_fd_sc_hd__nand2_1 _11435_ (.A(_05342_),
    .B(_05344_),
    .Y(_05623_));
 sky130_fd_sc_hd__a21bo_1 _11436_ (.A1(_05331_),
    .A2(_05333_),
    .B1_N(_05332_),
    .X(_05624_));
 sky130_fd_sc_hd__a22o_1 _11437_ (.A1(net626),
    .A2(net720),
    .B1(\dpath.alu.adder.in1[25] ),
    .B2(net630),
    .X(_05625_));
 sky130_fd_sc_hd__nand4_1 _11438_ (.A(net630),
    .B(net626),
    .C(net720),
    .D(\dpath.alu.adder.in1[25] ),
    .Y(_05626_));
 sky130_fd_sc_hd__nand4_2 _11439_ (.A(net622),
    .B(net721),
    .C(_05625_),
    .D(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__a22o_1 _11440_ (.A1(net622),
    .A2(net721),
    .B1(_05625_),
    .B2(_05626_),
    .X(_05628_));
 sky130_fd_sc_hd__nand3_1 _11441_ (.A(_05624_),
    .B(_05627_),
    .C(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__a21o_1 _11442_ (.A1(_05627_),
    .A2(_05628_),
    .B1(_05624_),
    .X(_05630_));
 sky130_fd_sc_hd__and3_1 _11443_ (.A(_05623_),
    .B(_05629_),
    .C(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__a21oi_1 _11444_ (.A1(_05629_),
    .A2(_05630_),
    .B1(_05623_),
    .Y(_05632_));
 sky130_fd_sc_hd__or4_2 _11445_ (.A(_05621_),
    .B(_05622_),
    .C(_05631_),
    .D(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__o22ai_2 _11446_ (.A1(_05621_),
    .A2(_05622_),
    .B1(_05631_),
    .B2(_05632_),
    .Y(_05634_));
 sky130_fd_sc_hd__nand3_1 _11447_ (.A(_05349_),
    .B(_05633_),
    .C(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__a21o_1 _11448_ (.A1(_05633_),
    .A2(_05634_),
    .B1(_05349_),
    .X(_05636_));
 sky130_fd_sc_hd__or4bb_2 _11449_ (.A(_05610_),
    .B(_05611_),
    .C_N(_05635_),
    .D_N(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__a2bb2o_1 _11450_ (.A1_N(_05610_),
    .A2_N(_05611_),
    .B1(_05635_),
    .B2(_05636_),
    .X(_05638_));
 sky130_fd_sc_hd__o211ai_2 _11451_ (.A1(_05351_),
    .A2(_05372_),
    .B1(_05637_),
    .C1(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a211o_1 _11452_ (.A1(_05637_),
    .A2(_05638_),
    .B1(_05351_),
    .C1(_05372_),
    .X(_05640_));
 sky130_fd_sc_hd__nand2_1 _11453_ (.A(_05639_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__xnor2_1 _11454_ (.A(_05592_),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__nor2_1 _11455_ (.A(_05375_),
    .B(_05409_),
    .Y(_05643_));
 sky130_fd_sc_hd__nand2b_1 _11456_ (.A_N(_05643_),
    .B(_05642_),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _11457_ (.A(_05642_),
    .B(_05643_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2b_1 _11458_ (.A_N(_05557_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__xor2_1 _11459_ (.A(_05557_),
    .B(_05645_),
    .X(_05647_));
 sky130_fd_sc_hd__nor2_1 _11460_ (.A(_05411_),
    .B(_05453_),
    .Y(_05648_));
 sky130_fd_sc_hd__xor2_1 _11461_ (.A(_05647_),
    .B(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__nand2b_1 _11462_ (.A_N(_05516_),
    .B(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__xnor2_1 _11463_ (.A(_05516_),
    .B(_05649_),
    .Y(_05651_));
 sky130_fd_sc_hd__o21a_1 _11464_ (.A1(_05455_),
    .A2(_05458_),
    .B1(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__nor3_1 _11465_ (.A(_05455_),
    .B(_05458_),
    .C(_05651_),
    .Y(_05653_));
 sky130_fd_sc_hd__nor2_1 _11466_ (.A(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__xor2_2 _11467_ (.A(_05515_),
    .B(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__or2_1 _11468_ (.A(_05461_),
    .B(_05463_),
    .X(_05656_));
 sky130_fd_sc_hd__nand2b_1 _11469_ (.A_N(_05655_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__xnor2_2 _11470_ (.A(_05655_),
    .B(_05656_),
    .Y(_05658_));
 sky130_fd_sc_hd__or2_1 _11471_ (.A(_05514_),
    .B(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__o311ai_4 _11472_ (.A1(_05287_),
    .A2(_05290_),
    .A3(_05466_),
    .B1(_05468_),
    .C1(_05658_),
    .Y(_05660_));
 sky130_fd_sc_hd__and3_1 _11473_ (.A(_02239_),
    .B(_05659_),
    .C(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__a221o_1 _11474_ (.A1(net3336),
    .A2(net486),
    .B1(_05512_),
    .B2(_05513_),
    .C1(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__a21oi_4 _11475_ (.A1(_02095_),
    .A2(net3337),
    .B1(_05510_),
    .Y(_05663_));
 sky130_fd_sc_hd__nor2_1 _11476_ (.A(net374),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _11477_ (.A(net578),
    .B(net3283),
    .Y(_05665_));
 sky130_fd_sc_hd__or2_1 _11478_ (.A(net578),
    .B(net3283),
    .X(_05666_));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_05665_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__a211o_1 _11480_ (.A1(_05298_),
    .A2(_05300_),
    .B1(_05479_),
    .C1(_05297_),
    .X(_05668_));
 sky130_fd_sc_hd__and2_1 _11481_ (.A(_05296_),
    .B(_05480_),
    .X(_05669_));
 sky130_fd_sc_hd__nand2_1 _11482_ (.A(_05668_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__a21o_1 _11483_ (.A1(_05668_),
    .A2(_05669_),
    .B1(_05667_),
    .X(_05671_));
 sky130_fd_sc_hd__xor2_1 _11484_ (.A(_05667_),
    .B(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__nor2_1 _11485_ (.A(net366),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__nand2_1 _11486_ (.A(net251),
    .B(_05484_),
    .Y(_05674_));
 sky130_fd_sc_hd__o211a_1 _11487_ (.A1(net251),
    .A2(_05484_),
    .B1(_05674_),
    .C1(net362),
    .X(_05675_));
 sky130_fd_sc_hd__a2111o_1 _11488_ (.A1(net3223),
    .A2(net404),
    .B1(net454),
    .C1(_05673_),
    .D1(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__o221a_1 _11489_ (.A1(net251),
    .A2(net446),
    .B1(_05664_),
    .B2(net3224),
    .C1(net858),
    .X(_00666_));
 sky130_fd_sc_hd__a21oi_1 _11490_ (.A1(net3246),
    .A2(_05674_),
    .B1(_01958_),
    .Y(_05677_));
 sky130_fd_sc_hd__o21a_1 _11491_ (.A1(net3246),
    .A2(_05674_),
    .B1(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__mux4_1 _11492_ (.A0(\dpath.RF.R[16][31] ),
    .A1(\dpath.RF.R[17][31] ),
    .A2(\dpath.RF.R[18][31] ),
    .A3(\dpath.RF.R[19][31] ),
    .S0(net575),
    .S1(net556),
    .X(_05679_));
 sky130_fd_sc_hd__nor2_1 _11493_ (.A(net536),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__mux4_1 _11494_ (.A0(\dpath.RF.R[20][31] ),
    .A1(\dpath.RF.R[21][31] ),
    .A2(\dpath.RF.R[22][31] ),
    .A3(\dpath.RF.R[23][31] ),
    .S0(net574),
    .S1(net555),
    .X(_05681_));
 sky130_fd_sc_hd__nor2_1 _11495_ (.A(net516),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__mux4_1 _11496_ (.A0(\dpath.RF.R[28][31] ),
    .A1(\dpath.RF.R[29][31] ),
    .A2(\dpath.RF.R[30][31] ),
    .A3(\dpath.RF.R[31][31] ),
    .S0(net575),
    .S1(net556),
    .X(_05683_));
 sky130_fd_sc_hd__nor2_1 _11497_ (.A(net516),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__mux4_1 _11498_ (.A0(\dpath.RF.R[24][31] ),
    .A1(\dpath.RF.R[25][31] ),
    .A2(\dpath.RF.R[26][31] ),
    .A3(\dpath.RF.R[27][31] ),
    .S0(net574),
    .S1(net555),
    .X(_05685_));
 sky130_fd_sc_hd__o21ai_1 _11499_ (.A1(net536),
    .A2(_05685_),
    .B1(net527),
    .Y(_05686_));
 sky130_fd_sc_hd__o32a_1 _11500_ (.A1(net526),
    .A2(_05680_),
    .A3(_05682_),
    .B1(_05684_),
    .B2(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__mux4_1 _11501_ (.A0(\dpath.RF.R[0][31] ),
    .A1(\dpath.RF.R[1][31] ),
    .A2(\dpath.RF.R[2][31] ),
    .A3(\dpath.RF.R[3][31] ),
    .S0(net575),
    .S1(net556),
    .X(_05688_));
 sky130_fd_sc_hd__nor2_1 _11502_ (.A(net537),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__mux4_1 _11503_ (.A0(\dpath.RF.R[4][31] ),
    .A1(\dpath.RF.R[5][31] ),
    .A2(\dpath.RF.R[6][31] ),
    .A3(\dpath.RF.R[7][31] ),
    .S0(net574),
    .S1(net555),
    .X(_05690_));
 sky130_fd_sc_hd__nor2_1 _11504_ (.A(net515),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__mux4_1 _11505_ (.A0(\dpath.RF.R[12][31] ),
    .A1(\dpath.RF.R[13][31] ),
    .A2(\dpath.RF.R[14][31] ),
    .A3(\dpath.RF.R[15][31] ),
    .S0(net574),
    .S1(net555),
    .X(_05692_));
 sky130_fd_sc_hd__mux4_1 _11506_ (.A0(\dpath.RF.R[8][31] ),
    .A1(\dpath.RF.R[9][31] ),
    .A2(\dpath.RF.R[10][31] ),
    .A3(\dpath.RF.R[11][31] ),
    .S0(net574),
    .S1(net555),
    .X(_05693_));
 sky130_fd_sc_hd__or2_1 _11507_ (.A(net537),
    .B(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__o211a_1 _11508_ (.A1(net515),
    .A2(_05692_),
    .B1(_05694_),
    .C1(net526),
    .X(_05695_));
 sky130_fd_sc_hd__nor2_1 _11509_ (.A(net520),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__o31a_1 _11510_ (.A1(net526),
    .A2(_05689_),
    .A3(_05691_),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__a211o_1 _11511_ (.A1(net520),
    .A2(_05687_),
    .B1(_05697_),
    .C1(net483),
    .X(_05698_));
 sky130_fd_sc_hd__nor2_1 _11512_ (.A(net372),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__mux2_2 _11513_ (.A0(net3664),
    .A1(net25),
    .S(net480),
    .X(_05700_));
 sky130_fd_sc_hd__a221o_1 _11514_ (.A1(net655),
    .A2(net369),
    .B1(net367),
    .B2(_05700_),
    .C1(_05699_),
    .X(_05701_));
 sky130_fd_sc_hd__a21oi_1 _11515_ (.A1(_01882_),
    .A2(_05512_),
    .B1(_01907_),
    .Y(_05702_));
 sky130_fd_sc_hd__a31o_1 _11516_ (.A1(_01882_),
    .A2(_01907_),
    .A3(_05512_),
    .B1(net469),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_1 _11517_ (.A(net768),
    .B(\dpath.alu.adder.in0[26] ),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_1 _11518_ (.A(_05542_),
    .B(_05544_),
    .Y(_05705_));
 sky130_fd_sc_hd__a21oi_1 _11519_ (.A1(_05569_),
    .A2(_05570_),
    .B1(_05572_),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ba_1 _11520_ (.A1(_05515_),
    .A2(_05653_),
    .B1_N(_05652_),
    .X(_05707_));
 sky130_fd_sc_hd__xnor2_1 _11521_ (.A(_05706_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__xnor2_1 _11522_ (.A(_05705_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__xnor2_1 _11523_ (.A(_05704_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__nor2_1 _11524_ (.A(_05546_),
    .B(_05548_),
    .Y(_05711_));
 sky130_fd_sc_hd__o21a_1 _11525_ (.A1(_05647_),
    .A2(_05648_),
    .B1(_05650_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _11526_ (.A(net777),
    .B(\dpath.alu.adder.in0[28] ),
    .Y(_05713_));
 sky130_fd_sc_hd__xor2_1 _11527_ (.A(_05712_),
    .B(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__xnor2_1 _11528_ (.A(_05711_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__xnor2_1 _11529_ (.A(_05710_),
    .B(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__o211ai_1 _11530_ (.A1(_05554_),
    .A2(_05556_),
    .B1(net784),
    .C1(\dpath.alu.adder.in0[30] ),
    .Y(_05717_));
 sky130_fd_sc_hd__a211o_1 _11531_ (.A1(net784),
    .A2(\dpath.alu.adder.in0[30] ),
    .B1(_05554_),
    .C1(_05556_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2_1 _11532_ (.A(_05717_),
    .B(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__o21ba_1 _11533_ (.A1(_05534_),
    .A2(_05551_),
    .B1_N(_05550_),
    .X(_05720_));
 sky130_fd_sc_hd__o21ba_1 _11534_ (.A1(_05527_),
    .A2(_05528_),
    .B1_N(_05526_),
    .X(_05721_));
 sky130_fd_sc_hd__xnor2_1 _11535_ (.A(_05720_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__nand2_1 _11536_ (.A(net739),
    .B(net588),
    .Y(_05723_));
 sky130_fd_sc_hd__nand2_1 _11537_ (.A(net735),
    .B(net592),
    .Y(_05724_));
 sky130_fd_sc_hd__xnor2_1 _11538_ (.A(_05723_),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__xnor2_1 _11539_ (.A(_05722_),
    .B(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__xnor2_1 _11540_ (.A(_05719_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2_1 _11541_ (.A(net764),
    .B(\dpath.alu.adder.in0[25] ),
    .Y(_05728_));
 sky130_fd_sc_hd__nand2_1 _11542_ (.A(net743),
    .B(net585),
    .Y(_05729_));
 sky130_fd_sc_hd__a211oi_1 _11543_ (.A1(net738),
    .A2(net590),
    .B1(_05608_),
    .C1(_05610_),
    .Y(_05730_));
 sky130_fd_sc_hd__o211a_1 _11544_ (.A1(_05608_),
    .A2(_05610_),
    .B1(net738),
    .C1(net589),
    .X(_05731_));
 sky130_fd_sc_hd__nor2_1 _11545_ (.A(_05730_),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__xnor2_1 _11546_ (.A(_05729_),
    .B(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__xnor2_1 _11547_ (.A(_05728_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__xnor2_1 _11548_ (.A(_05727_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__o31ai_1 _11549_ (.A1(_05559_),
    .A2(_05587_),
    .A3(_05588_),
    .B1(_05591_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand2_1 _11550_ (.A(net772),
    .B(\dpath.alu.adder.in0[27] ),
    .Y(_05737_));
 sky130_fd_sc_hd__nand2_1 _11551_ (.A(_05604_),
    .B(_05606_),
    .Y(_05738_));
 sky130_fd_sc_hd__xor2_1 _11552_ (.A(_05737_),
    .B(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__xnor2_1 _11553_ (.A(_05736_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__xnor2_1 _11554_ (.A(_05735_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__xnor2_1 _11555_ (.A(_05716_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__a31o_1 _11556_ (.A1(net759),
    .A2(net580),
    .A3(_05562_),
    .B1(_05561_),
    .X(_05743_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_05644_),
    .B(_05646_),
    .Y(_05744_));
 sky130_fd_sc_hd__xnor2_1 _11558_ (.A(_05743_),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__a31o_1 _11559_ (.A1(net780),
    .A2(\dpath.alu.adder.in0[28] ),
    .A3(_05522_),
    .B1(_05521_),
    .X(_05746_));
 sky130_fd_sc_hd__a21bo_1 _11560_ (.A1(\dpath.alu.adder.in1[6] ),
    .A2(net579),
    .B1_N(_05540_),
    .X(_05747_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(net763),
    .B(\dpath.alu.adder.in0[24] ),
    .Y(_05748_));
 sky130_fd_sc_hd__mux2_1 _11562_ (.A0(_05747_),
    .A1(_05540_),
    .S(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__nand2_1 _11563_ (.A(net614),
    .B(net722),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_1 _11564_ (.A(net747),
    .B(net583),
    .Y(_05751_));
 sky130_fd_sc_hd__xor2_1 _11565_ (.A(_05750_),
    .B(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__nand2_1 _11566_ (.A(net780),
    .B(\dpath.alu.adder.in0[29] ),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(net787),
    .B(\dpath.alu.adder.in0[31] ),
    .Y(_05754_));
 sky130_fd_sc_hd__xor2_1 _11568_ (.A(_05753_),
    .B(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__nand2_1 _11569_ (.A(net610),
    .B(net723),
    .Y(_05756_));
 sky130_fd_sc_hd__nand2_1 _11570_ (.A(net605),
    .B(net726),
    .Y(_05757_));
 sky130_fd_sc_hd__a31o_1 _11571_ (.A1(_05624_),
    .A2(_05627_),
    .A3(_05628_),
    .B1(_05631_),
    .X(_05758_));
 sky130_fd_sc_hd__xnor2_1 _11572_ (.A(_05757_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__nand2_1 _11573_ (.A(net622),
    .B(net720),
    .Y(_05760_));
 sky130_fd_sc_hd__nand2_1 _11574_ (.A(_05613_),
    .B(_05615_),
    .Y(_05761_));
 sky130_fd_sc_hd__xnor2_1 _11575_ (.A(_05619_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__xnor2_1 _11576_ (.A(_05760_),
    .B(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2_1 _11577_ (.A(net644),
    .B(\dpath.alu.adder.in1[29] ),
    .Y(_05764_));
 sky130_fd_sc_hd__and3_1 _11578_ (.A(net648),
    .B(\dpath.alu.adder.in1[30] ),
    .C(_05330_),
    .X(_05765_));
 sky130_fd_sc_hd__xnor2_1 _11579_ (.A(_05764_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__nand2_1 _11580_ (.A(net652),
    .B(\dpath.alu.adder.in1[31] ),
    .Y(_05767_));
 sky130_fd_sc_hd__xnor2_1 _11581_ (.A(_05766_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__xnor2_1 _11582_ (.A(_05763_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__xnor2_1 _11583_ (.A(_05759_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__xnor2_1 _11584_ (.A(_05756_),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_2 _11585_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05566_),
    .Y(_05772_));
 sky130_fd_sc_hd__nand2_1 _11586_ (.A(net756),
    .B(net580),
    .Y(_05773_));
 sky130_fd_sc_hd__xnor2_2 _11587_ (.A(_05772_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(net599),
    .B(net730),
    .Y(_05775_));
 sky130_fd_sc_hd__a21bo_1 _11589_ (.A1(net630),
    .A2(net720),
    .B1_N(_05627_),
    .X(_05776_));
 sky130_fd_sc_hd__nand2_1 _11590_ (.A(net626),
    .B(\dpath.alu.adder.in1[25] ),
    .Y(_05777_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(_05776_),
    .A1(_05627_),
    .S(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__xor2_1 _11592_ (.A(_05775_),
    .B(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__nand2b_1 _11593_ (.A_N(_05622_),
    .B(_05633_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand2_1 _11594_ (.A(net618),
    .B(net721),
    .Y(_05781_));
 sky130_fd_sc_hd__xor2_1 _11595_ (.A(_05780_),
    .B(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__nand2_1 _11596_ (.A(net640),
    .B(\dpath.alu.adder.in1[28] ),
    .Y(_05783_));
 sky130_fd_sc_hd__nand2_1 _11597_ (.A(net634),
    .B(\dpath.alu.adder.in1[27] ),
    .Y(_05784_));
 sky130_fd_sc_hd__nand2_1 _11598_ (.A(net630),
    .B(\dpath.alu.adder.in1[26] ),
    .Y(_05785_));
 sky130_fd_sc_hd__xnor2_1 _11599_ (.A(_05784_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__xnor2_1 _11600_ (.A(_05783_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__xnor2_1 _11601_ (.A(_05782_),
    .B(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__xnor2_1 _11602_ (.A(_05779_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__xnor2_1 _11603_ (.A(_05774_),
    .B(_05789_),
    .Y(_05790_));
 sky130_fd_sc_hd__xnor2_1 _11604_ (.A(_05771_),
    .B(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _11605_ (.A(net607),
    .B(net725),
    .Y(_05792_));
 sky130_fd_sc_hd__nand2_1 _11606_ (.A(net601),
    .B(net728),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_1 _11607_ (.A(_05635_),
    .B(_05637_),
    .Y(_05794_));
 sky130_fd_sc_hd__nand2_1 _11608_ (.A(_05600_),
    .B(_05602_),
    .Y(_05795_));
 sky130_fd_sc_hd__xor2_1 _11609_ (.A(_05794_),
    .B(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__xnor2_1 _11610_ (.A(_05793_),
    .B(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__xnor2_1 _11611_ (.A(_05792_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__xnor2_2 _11612_ (.A(_05791_),
    .B(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__xnor2_1 _11613_ (.A(_05755_),
    .B(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__nand2_1 _11614_ (.A(net753),
    .B(net581),
    .Y(_05801_));
 sky130_fd_sc_hd__a31o_1 _11615_ (.A1(net787),
    .A2(\dpath.alu.adder.in0[30] ),
    .A3(_05532_),
    .B1(_05530_),
    .X(_05802_));
 sky130_fd_sc_hd__a31o_1 _11616_ (.A1(_05582_),
    .A2(_05583_),
    .A3(_05584_),
    .B1(_05587_),
    .X(_05803_));
 sky130_fd_sc_hd__xnor2_1 _11617_ (.A(_05802_),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__xnor2_1 _11618_ (.A(_05801_),
    .B(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__a21boi_1 _11619_ (.A1(_05592_),
    .A2(_05640_),
    .B1_N(_05639_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _11620_ (.A(net759),
    .B(net579),
    .Y(_05807_));
 sky130_fd_sc_hd__xor2_1 _11621_ (.A(_05806_),
    .B(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__a21bo_1 _11622_ (.A1(net599),
    .A2(net735),
    .B1_N(_05578_),
    .X(_05809_));
 sky130_fd_sc_hd__nand2_1 _11623_ (.A(net595),
    .B(net733),
    .Y(_05810_));
 sky130_fd_sc_hd__mux2_1 _11624_ (.A0(_05809_),
    .A1(_05578_),
    .S(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__a31o_1 _11625_ (.A1(net602),
    .A2(net730),
    .A3(_05596_),
    .B1(_05595_),
    .X(_05812_));
 sky130_fd_sc_hd__and3_1 _11626_ (.A(_05580_),
    .B(_05582_),
    .C(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__a21oi_1 _11627_ (.A1(_05580_),
    .A2(_05582_),
    .B1(_05812_),
    .Y(_05814_));
 sky130_fd_sc_hd__or2_1 _11628_ (.A(_05813_),
    .B(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__xnor2_1 _11629_ (.A(_05811_),
    .B(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__xnor2_1 _11630_ (.A(_05808_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__xnor2_1 _11631_ (.A(_05805_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__xnor2_1 _11632_ (.A(_05800_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__xnor2_1 _11633_ (.A(_05752_),
    .B(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__xnor2_1 _11634_ (.A(_05749_),
    .B(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__xnor2_1 _11635_ (.A(_05746_),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__xnor2_1 _11636_ (.A(_05745_),
    .B(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__xnor2_2 _11637_ (.A(_05742_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__a21oi_1 _11638_ (.A1(_05657_),
    .A2(_05660_),
    .B1(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__a311o_1 _11639_ (.A1(_05657_),
    .A2(_05660_),
    .A3(_05824_),
    .B1(_05825_),
    .C1(net485),
    .X(_05826_));
 sky130_fd_sc_hd__o21a_1 _11640_ (.A1(net3679),
    .A2(_02071_),
    .B1(net469),
    .X(_05827_));
 sky130_fd_sc_hd__a2bb2o_2 _11641_ (.A1_N(_05702_),
    .A2_N(_05703_),
    .B1(_05826_),
    .B2(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__a21oi_4 _11642_ (.A1(_02095_),
    .A2(_05828_),
    .B1(_05701_),
    .Y(_05829_));
 sky130_fd_sc_hd__nand2_1 _11643_ (.A(net3422),
    .B(_01952_),
    .Y(_05830_));
 sky130_fd_sc_hd__nor2_1 _11644_ (.A(net578),
    .B(net3184),
    .Y(_05831_));
 sky130_fd_sc_hd__and2_1 _11645_ (.A(net578),
    .B(net3184),
    .X(_05832_));
 sky130_fd_sc_hd__o211a_1 _11646_ (.A1(_05831_),
    .A2(_05832_),
    .B1(_05665_),
    .C1(_05671_),
    .X(_05833_));
 sky130_fd_sc_hd__a211oi_1 _11647_ (.A1(_05665_),
    .A2(_05671_),
    .B1(_05831_),
    .C1(_05832_),
    .Y(_05834_));
 sky130_fd_sc_hd__o32a_1 _11648_ (.A1(net366),
    .A2(_05833_),
    .A3(_05834_),
    .B1(_05829_),
    .B2(net374),
    .X(_05835_));
 sky130_fd_sc_hd__a31o_1 _11649_ (.A1(_01958_),
    .A2(_05830_),
    .A3(_05835_),
    .B1(_05678_),
    .X(_05836_));
 sky130_fd_sc_hd__nor2_1 _11650_ (.A(net3246),
    .B(net446),
    .Y(_05837_));
 sky130_fd_sc_hd__a211oi_1 _11651_ (.A1(net446),
    .A2(net3423),
    .B1(_05837_),
    .C1(net880),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_4 _11652_ (.A(_01820_),
    .B(_02014_),
    .Y(_05838_));
 sky130_fd_sc_hd__mux2_1 _11653_ (.A0(net719),
    .A1(net2096),
    .S(net389),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(net716),
    .A1(net3068),
    .S(net389),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _11655_ (.A0(net715),
    .A1(net3146),
    .S(net389),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _11656_ (.A0(net713),
    .A1(net2876),
    .S(net389),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _11657_ (.A0(net711),
    .A1(net2526),
    .S(net389),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(net709),
    .A1(net2036),
    .S(net389),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _11659_ (.A0(net707),
    .A1(net3136),
    .S(net389),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(net705),
    .A1(net2854),
    .S(net389),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(net702),
    .A1(net2462),
    .S(net389),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(net701),
    .A1(net3004),
    .S(net389),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(net699),
    .A1(net2118),
    .S(net389),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(net696),
    .A1(net3154),
    .S(net389),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _11665_ (.A0(net695),
    .A1(net2698),
    .S(net389),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _11666_ (.A0(net692),
    .A1(net1964),
    .S(net389),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(net691),
    .A1(net2450),
    .S(net389),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(\dpath.RF.wdata[15] ),
    .A1(net2052),
    .S(net389),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _11669_ (.A0(net687),
    .A1(net2518),
    .S(net390),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(net685),
    .A1(net1768),
    .S(net390),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _11671_ (.A0(net683),
    .A1(net1482),
    .S(net390),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(net681),
    .A1(net2460),
    .S(net390),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _11673_ (.A0(net679),
    .A1(net2658),
    .S(net390),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(net676),
    .A1(net2672),
    .S(net390),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _11675_ (.A0(net3714),
    .A1(net1624),
    .S(net390),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _11676_ (.A0(net672),
    .A1(net3066),
    .S(net390),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _11677_ (.A0(net670),
    .A1(net2822),
    .S(net390),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(net667),
    .A1(net2490),
    .S(net390),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(net664),
    .A1(net3196),
    .S(net390),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(net663),
    .A1(net2408),
    .S(net390),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(net660),
    .A1(net1894),
    .S(net390),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _11682_ (.A0(net659),
    .A1(net2082),
    .S(net390),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(net656),
    .A1(net2288),
    .S(net390),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(net655),
    .A1(net2166),
    .S(net390),
    .X(_00699_));
 sky130_fd_sc_hd__or2_1 _11685_ (.A(net45),
    .B(net453),
    .X(_05839_));
 sky130_fd_sc_hd__o211a_1 _11686_ (.A1(net3432),
    .A2(net446),
    .B1(_05839_),
    .C1(net854),
    .X(_00700_));
 sky130_fd_sc_hd__or2_1 _11687_ (.A(net46),
    .B(net453),
    .X(_05840_));
 sky130_fd_sc_hd__o211a_1 _11688_ (.A1(net3393),
    .A2(net448),
    .B1(_05840_),
    .C1(net854),
    .X(_00701_));
 sky130_fd_sc_hd__or2_1 _11689_ (.A(net47),
    .B(net453),
    .X(_05841_));
 sky130_fd_sc_hd__o211a_1 _11690_ (.A1(net3403),
    .A2(net448),
    .B1(_05841_),
    .C1(net854),
    .X(_00702_));
 sky130_fd_sc_hd__or2_1 _11691_ (.A(net48),
    .B(net453),
    .X(_05842_));
 sky130_fd_sc_hd__o211a_1 _11692_ (.A1(net3285),
    .A2(net448),
    .B1(_05842_),
    .C1(net856),
    .X(_00703_));
 sky130_fd_sc_hd__or2_1 _11693_ (.A(net49),
    .B(net453),
    .X(_05843_));
 sky130_fd_sc_hd__o211a_1 _11694_ (.A1(net3349),
    .A2(net448),
    .B1(_05843_),
    .C1(net856),
    .X(_00704_));
 sky130_fd_sc_hd__or3_4 _11695_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(_01779_),
    .C(\ctrl.c2d_rf_waddr_W[4] ),
    .X(_05844_));
 sky130_fd_sc_hd__nor2_4 _11696_ (.A(_01830_),
    .B(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__mux2_1 _11697_ (.A0(net1184),
    .A1(net718),
    .S(net387),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(net2962),
    .A1(net717),
    .S(net387),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _11699_ (.A0(net2648),
    .A1(net714),
    .S(net387),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(net1834),
    .A1(net712),
    .S(net387),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _11701_ (.A0(net1378),
    .A1(net710),
    .S(net387),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(net1684),
    .A1(net708),
    .S(net387),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _11703_ (.A0(net2736),
    .A1(net706),
    .S(net387),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(net2918),
    .A1(net704),
    .S(net387),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _11705_ (.A0(net1604),
    .A1(net703),
    .S(net387),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(net2994),
    .A1(net700),
    .S(net387),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(net2270),
    .A1(net698),
    .S(net387),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(net2546),
    .A1(net697),
    .S(net387),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _11709_ (.A0(net1904),
    .A1(net694),
    .S(net387),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _11710_ (.A0(net1620),
    .A1(net693),
    .S(net387),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(net2100),
    .A1(net690),
    .S(net387),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _11712_ (.A0(net1564),
    .A1(net688),
    .S(net387),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _11713_ (.A0(net2308),
    .A1(net686),
    .S(net388),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(net2666),
    .A1(net684),
    .S(net388),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _11715_ (.A0(net2342),
    .A1(net682),
    .S(net388),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _11716_ (.A0(net1444),
    .A1(net680),
    .S(net388),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _11717_ (.A0(net3002),
    .A1(net677),
    .S(net388),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(net2378),
    .A1(net675),
    .S(net388),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(net2120),
    .A1(net673),
    .S(net388),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(net1544),
    .A1(net671),
    .S(net388),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(net2806),
    .A1(net668),
    .S(net388),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _11722_ (.A0(net1326),
    .A1(net666),
    .S(net388),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _11723_ (.A0(net1578),
    .A1(net665),
    .S(net388),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _11724_ (.A0(net1744),
    .A1(\dpath.RF.wdata[27] ),
    .S(net388),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(net1244),
    .A1(net661),
    .S(net388),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(net1308),
    .A1(net658),
    .S(net388),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _11727_ (.A0(net1770),
    .A1(net657),
    .S(net388),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _11728_ (.A0(net1280),
    .A1(\dpath.RF.wdata[31] ),
    .S(net388),
    .X(_00736_));
 sky130_fd_sc_hd__or3_4 _11729_ (.A(\ctrl.c2d_rf_waddr_W[2] ),
    .B(_01779_),
    .C(_01780_),
    .X(_05846_));
 sky130_fd_sc_hd__or2_4 _11730_ (.A(_01830_),
    .B(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__mux2_1 _11731_ (.A0(\dpath.RF.wdata[0] ),
    .A1(net1334),
    .S(net386),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(net716),
    .A1(net2884),
    .S(net386),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _11733_ (.A0(net1374),
    .A1(net3708),
    .S(net386),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(net713),
    .A1(net3058),
    .S(net386),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(net711),
    .A1(net3090),
    .S(net386),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(net709),
    .A1(net3134),
    .S(net386),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _11737_ (.A0(net706),
    .A1(net2902),
    .S(net386),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(net705),
    .A1(net1796),
    .S(net386),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _11739_ (.A0(net702),
    .A1(net2680),
    .S(net386),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(net701),
    .A1(net1644),
    .S(net386),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(net699),
    .A1(net2878),
    .S(net386),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(net696),
    .A1(net3072),
    .S(net386),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _11743_ (.A0(net695),
    .A1(net3160),
    .S(net386),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _11744_ (.A0(net692),
    .A1(net2396),
    .S(net386),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(net691),
    .A1(net1548),
    .S(net386),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(net689),
    .A1(net2468),
    .S(net385),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(net687),
    .A1(net2818),
    .S(net385),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(net685),
    .A1(net1588),
    .S(net385),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(net683),
    .A1(net1962),
    .S(net385),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(net681),
    .A1(net2528),
    .S(net385),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _11751_ (.A0(net679),
    .A1(net2356),
    .S(net385),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(net676),
    .A1(net2306),
    .S(net385),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(net674),
    .A1(net2772),
    .S(net385),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(net672),
    .A1(net2382),
    .S(net385),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(net670),
    .A1(net2044),
    .S(net385),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _11756_ (.A0(net667),
    .A1(net1878),
    .S(net385),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(net664),
    .A1(net1722),
    .S(net385),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(net663),
    .A1(net1764),
    .S(net385),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _11759_ (.A0(net660),
    .A1(net2386),
    .S(net385),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(net659),
    .A1(net3094),
    .S(net385),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _11761_ (.A0(net656),
    .A1(net2790),
    .S(net385),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(net655),
    .A1(net2536),
    .S(_05847_),
    .X(_00768_));
 sky130_fd_sc_hd__nor2_4 _11763_ (.A(_01823_),
    .B(_01832_),
    .Y(_05848_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(net2786),
    .A1(net718),
    .S(net431),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _11765_ (.A0(net1802),
    .A1(net717),
    .S(net431),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(net2296),
    .A1(net714),
    .S(net431),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(net1866),
    .A1(net712),
    .S(net431),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(net1756),
    .A1(net710),
    .S(net431),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(net2236),
    .A1(net708),
    .S(net431),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(net2844),
    .A1(net706),
    .S(net431),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(net2440),
    .A1(net705),
    .S(net431),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(net2212),
    .A1(net702),
    .S(net431),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _11773_ (.A0(net2474),
    .A1(net700),
    .S(net431),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _11774_ (.A0(net2086),
    .A1(net698),
    .S(net431),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _11775_ (.A0(net2084),
    .A1(net697),
    .S(net431),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _11776_ (.A0(net2090),
    .A1(net694),
    .S(net431),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _11777_ (.A0(net1592),
    .A1(net693),
    .S(net431),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _11778_ (.A0(net2484),
    .A1(net690),
    .S(net431),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _11779_ (.A0(net2332),
    .A1(net688),
    .S(net431),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(net1480),
    .A1(net686),
    .S(net432),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _11781_ (.A0(net2292),
    .A1(net684),
    .S(net432),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _11782_ (.A0(net1436),
    .A1(net682),
    .S(net432),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _11783_ (.A0(net1508),
    .A1(net681),
    .S(net432),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(net2804),
    .A1(net677),
    .S(net432),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _11785_ (.A0(net2400),
    .A1(net676),
    .S(net432),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _11786_ (.A0(net1402),
    .A1(net673),
    .S(net432),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _11787_ (.A0(net2018),
    .A1(net671),
    .S(net432),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _11788_ (.A0(net1206),
    .A1(net669),
    .S(net432),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _11789_ (.A0(net1380),
    .A1(net666),
    .S(net432),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(net2140),
    .A1(net665),
    .S(net432),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _11791_ (.A0(net1518),
    .A1(net663),
    .S(net432),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _11792_ (.A0(net1598),
    .A1(net661),
    .S(net432),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _11793_ (.A0(net1928),
    .A1(net659),
    .S(net432),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _11794_ (.A0(net1248),
    .A1(net657),
    .S(net432),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _11795_ (.A0(net1452),
    .A1(net654),
    .S(net432),
    .X(_00832_));
 sky130_fd_sc_hd__nor2_4 _11796_ (.A(_01823_),
    .B(_05844_),
    .Y(_05849_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(net1750),
    .A1(net718),
    .S(net429),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _11798_ (.A0(net2850),
    .A1(net717),
    .S(net429),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _11799_ (.A0(net1658),
    .A1(net714),
    .S(net429),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _11800_ (.A0(net1818),
    .A1(net712),
    .S(net429),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _11801_ (.A0(net1416),
    .A1(net710),
    .S(net429),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _11802_ (.A0(net2388),
    .A1(net708),
    .S(net429),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(net1890),
    .A1(net706),
    .S(net429),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _11804_ (.A0(net2410),
    .A1(net705),
    .S(net429),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _11805_ (.A0(net1270),
    .A1(net703),
    .S(net429),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _11806_ (.A0(net1464),
    .A1(net700),
    .S(net429),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(net1952),
    .A1(net698),
    .S(net429),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(net2592),
    .A1(net697),
    .S(net429),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(net2122),
    .A1(net694),
    .S(net429),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(net2046),
    .A1(net693),
    .S(net429),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(net1782),
    .A1(net690),
    .S(net429),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _11812_ (.A0(net2580),
    .A1(net688),
    .S(net429),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(net2278),
    .A1(net686),
    .S(net430),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _11814_ (.A0(net1246),
    .A1(net684),
    .S(net430),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(net2152),
    .A1(net682),
    .S(net430),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(net2452),
    .A1(net681),
    .S(net430),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(net1510),
    .A1(net677),
    .S(net430),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(net1218),
    .A1(\dpath.RF.wdata[21] ),
    .S(net430),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(net2960),
    .A1(net673),
    .S(net430),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(net1742),
    .A1(net671),
    .S(net430),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(net1814),
    .A1(net668),
    .S(net430),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(net1190),
    .A1(net666),
    .S(net430),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(net2704),
    .A1(net665),
    .S(net430),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _11824_ (.A0(net1376),
    .A1(net663),
    .S(net430),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(net1258),
    .A1(net661),
    .S(net430),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(net1622),
    .A1(net658),
    .S(net430),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(net1236),
    .A1(net657),
    .S(net430),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(net1682),
    .A1(net655),
    .S(net430),
    .X(_00864_));
 sky130_fd_sc_hd__nor2_4 _11829_ (.A(_01827_),
    .B(_02019_),
    .Y(_05850_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(net3084),
    .A1(net719),
    .S(net427),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(net1748),
    .A1(net3711),
    .S(net427),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(net1348),
    .A1(net715),
    .S(net427),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(net1852),
    .A1(net3271),
    .S(net427),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(net2512),
    .A1(net711),
    .S(net427),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _11835_ (.A0(net1330),
    .A1(net3678),
    .S(net427),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(net3710),
    .A1(net1360),
    .S(net427),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _11837_ (.A0(net1994),
    .A1(net704),
    .S(net427),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(net2682),
    .A1(net702),
    .S(net427),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _11839_ (.A0(net2198),
    .A1(\dpath.RF.wdata[9] ),
    .S(net427),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(net1860),
    .A1(net699),
    .S(net427),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _11841_ (.A0(net2144),
    .A1(net696),
    .S(net427),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(net1892),
    .A1(net695),
    .S(net427),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _11843_ (.A0(net1492),
    .A1(net692),
    .S(net427),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(net1686),
    .A1(net3716),
    .S(net427),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(net2142),
    .A1(net689),
    .S(net427),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(net2326),
    .A1(\dpath.RF.wdata[16] ),
    .S(net428),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _11847_ (.A0(net1954),
    .A1(net685),
    .S(net428),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(net2230),
    .A1(net683),
    .S(net428),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(net1616),
    .A1(net680),
    .S(net428),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(net2088),
    .A1(net678),
    .S(net428),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _11851_ (.A0(net1816),
    .A1(net675),
    .S(net428),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _11852_ (.A0(net1340),
    .A1(net674),
    .S(net428),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(net1502),
    .A1(net672),
    .S(net428),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(net1666),
    .A1(net668),
    .S(net428),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(net1972),
    .A1(net667),
    .S(net428),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(net2568),
    .A1(net664),
    .S(net428),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(net2668),
    .A1(net662),
    .S(net428),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(net1546),
    .A1(net660),
    .S(net428),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(net1772),
    .A1(net659),
    .S(net428),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _11860_ (.A0(net1382),
    .A1(net3712),
    .S(net428),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(net1364),
    .A1(net654),
    .S(net428),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_4 _11862_ (.A(_01823_),
    .B(_05846_),
    .Y(_05851_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(net2274),
    .A1(net719),
    .S(net426),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _11864_ (.A0(net1238),
    .A1(net716),
    .S(net426),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(net2148),
    .A1(net715),
    .S(net426),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _11866_ (.A0(net1614),
    .A1(net712),
    .S(net426),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(net1566),
    .A1(net710),
    .S(net426),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _11868_ (.A0(net2110),
    .A1(net709),
    .S(net426),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(net2184),
    .A1(net706),
    .S(net426),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _11870_ (.A0(net1438),
    .A1(net705),
    .S(net426),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(net1710),
    .A1(net702),
    .S(net426),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _11872_ (.A0(net1474),
    .A1(net701),
    .S(net426),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(net1324),
    .A1(net699),
    .S(net426),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(net2280),
    .A1(net696),
    .S(net426),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(net2810),
    .A1(net695),
    .S(net426),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(net2650),
    .A1(net692),
    .S(net426),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(net1910),
    .A1(net691),
    .S(net426),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(net1632),
    .A1(\dpath.RF.wdata[15] ),
    .S(net425),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _11879_ (.A0(net1882),
    .A1(net687),
    .S(net425),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(net2434),
    .A1(net685),
    .S(net425),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _11881_ (.A0(net1806),
    .A1(net683),
    .S(net425),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _11882_ (.A0(net1936),
    .A1(net681),
    .S(net425),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _11883_ (.A0(net1828),
    .A1(net679),
    .S(net425),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _11884_ (.A0(net2138),
    .A1(net676),
    .S(net425),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _11885_ (.A0(net1386),
    .A1(net674),
    .S(net425),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(net1220),
    .A1(\dpath.RF.wdata[23] ),
    .S(net425),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _11887_ (.A0(net2162),
    .A1(net670),
    .S(net425),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(net1226),
    .A1(net667),
    .S(net425),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _11889_ (.A0(net2428),
    .A1(net664),
    .S(net425),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(net1932),
    .A1(net663),
    .S(net425),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _11891_ (.A0(net1626),
    .A1(net660),
    .S(net425),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(net1408),
    .A1(net659),
    .S(net425),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _11893_ (.A0(net1550),
    .A1(net656),
    .S(net425),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _11894_ (.A0(net1466),
    .A1(net655),
    .S(_05851_),
    .X(_00928_));
 sky130_fd_sc_hd__or2_4 _11895_ (.A(_01821_),
    .B(_05844_),
    .X(_05852_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(net718),
    .A1(net2498),
    .S(net383),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _11897_ (.A0(net717),
    .A1(net3092),
    .S(net383),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(net714),
    .A1(net2912),
    .S(net383),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(net712),
    .A1(net3114),
    .S(net383),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(net710),
    .A1(net2294),
    .S(net383),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(net708),
    .A1(net2248),
    .S(net383),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _11902_ (.A0(net706),
    .A1(net2888),
    .S(net383),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _11903_ (.A0(net705),
    .A1(net2372),
    .S(net383),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(net703),
    .A1(net1946),
    .S(net383),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _11905_ (.A0(net700),
    .A1(net2480),
    .S(net383),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _11906_ (.A0(net698),
    .A1(net1862),
    .S(net383),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _11907_ (.A0(net697),
    .A1(net3158),
    .S(net383),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(net694),
    .A1(net2982),
    .S(net383),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _11909_ (.A0(net693),
    .A1(net2012),
    .S(net383),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(net690),
    .A1(net2530),
    .S(net383),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _11911_ (.A0(net688),
    .A1(net2302),
    .S(net383),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(net686),
    .A1(net3096),
    .S(net384),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(net684),
    .A1(net2812),
    .S(net384),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(net682),
    .A1(net2942),
    .S(net384),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(net681),
    .A1(net2846),
    .S(net384),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _11916_ (.A0(net677),
    .A1(net2632),
    .S(net384),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(\dpath.RF.wdata[21] ),
    .A1(net1760),
    .S(net384),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _11918_ (.A0(net673),
    .A1(net2956),
    .S(net384),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _11919_ (.A0(net671),
    .A1(net3024),
    .S(net384),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(net668),
    .A1(net2136),
    .S(net384),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(net666),
    .A1(net2792),
    .S(net384),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _11922_ (.A0(net665),
    .A1(net2798),
    .S(net384),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _11923_ (.A0(net662),
    .A1(net2000),
    .S(net384),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _11924_ (.A0(net661),
    .A1(net2904),
    .S(net384),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _11925_ (.A0(net658),
    .A1(net1982),
    .S(net384),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _11926_ (.A0(net657),
    .A1(net3164),
    .S(net384),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _11927_ (.A0(net655),
    .A1(net1886),
    .S(net384),
    .X(_00960_));
 sky130_fd_sc_hd__or2_4 _11928_ (.A(_01821_),
    .B(_05846_),
    .X(_05853_));
 sky130_fd_sc_hd__mux2_1 _11929_ (.A0(net718),
    .A1(net3148),
    .S(net382),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _11930_ (.A0(net716),
    .A1(net1900),
    .S(net382),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _11931_ (.A0(net715),
    .A1(net2074),
    .S(net382),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _11932_ (.A0(net712),
    .A1(net2204),
    .S(net382),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _11933_ (.A0(net710),
    .A1(net2776),
    .S(net382),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(net709),
    .A1(net2062),
    .S(net382),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _11935_ (.A0(net706),
    .A1(net2340),
    .S(net382),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(net705),
    .A1(net2690),
    .S(net382),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _11937_ (.A0(net702),
    .A1(net2032),
    .S(net382),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _11938_ (.A0(net701),
    .A1(net2416),
    .S(net382),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _11939_ (.A0(net1078),
    .A1(net3694),
    .S(net382),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(net696),
    .A1(net3022),
    .S(net382),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _11941_ (.A0(net695),
    .A1(net2856),
    .S(net382),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(net692),
    .A1(net3110),
    .S(net382),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(net691),
    .A1(net2192),
    .S(net382),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(net689),
    .A1(net2694),
    .S(net381),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _11945_ (.A0(net687),
    .A1(net2054),
    .S(net381),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _11946_ (.A0(net685),
    .A1(net2996),
    .S(net381),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(net683),
    .A1(net1758),
    .S(net381),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _11948_ (.A0(net681),
    .A1(net3162),
    .S(net381),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(net679),
    .A1(net2068),
    .S(net381),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _11950_ (.A0(net676),
    .A1(net2334),
    .S(net381),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(net674),
    .A1(net2258),
    .S(net381),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _11952_ (.A0(\dpath.RF.wdata[23] ),
    .A1(net2610),
    .S(net381),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(net670),
    .A1(net3142),
    .S(net381),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _11954_ (.A0(net667),
    .A1(net3054),
    .S(net381),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(net664),
    .A1(net2930),
    .S(net381),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _11956_ (.A0(net663),
    .A1(net1668),
    .S(net381),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _11957_ (.A0(net3704),
    .A1(net2524),
    .S(net381),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _11958_ (.A0(net659),
    .A1(net2112),
    .S(net381),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _11959_ (.A0(net656),
    .A1(net1690),
    .S(net381),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _11960_ (.A0(net655),
    .A1(net2284),
    .S(_05853_),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_4 _11961_ (.A(_02019_),
    .B(_05844_),
    .Y(_05854_));
 sky130_fd_sc_hd__mux2_1 _11962_ (.A0(net1484),
    .A1(net718),
    .S(net423),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(net2692),
    .A1(net717),
    .S(net423),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _11964_ (.A0(net2840),
    .A1(net714),
    .S(net423),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(net1998),
    .A1(net712),
    .S(net423),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _11966_ (.A0(net2470),
    .A1(net710),
    .S(net423),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(net2246),
    .A1(net708),
    .S(net423),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _11968_ (.A0(net1948),
    .A1(net706),
    .S(net423),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(net2834),
    .A1(net704),
    .S(net423),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(net2366),
    .A1(net703),
    .S(net423),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(net1560),
    .A1(net700),
    .S(net423),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _11972_ (.A0(net2478),
    .A1(net698),
    .S(net423),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(net2500),
    .A1(net697),
    .S(net423),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _11974_ (.A0(net2272),
    .A1(net694),
    .S(net423),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _11975_ (.A0(net1680),
    .A1(net693),
    .S(net423),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _11976_ (.A0(net1534),
    .A1(net690),
    .S(net423),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _11977_ (.A0(net1832),
    .A1(net688),
    .S(net423),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _11978_ (.A0(net2476),
    .A1(net686),
    .S(net424),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _11979_ (.A0(net2202),
    .A1(net684),
    .S(net424),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(net2006),
    .A1(net682),
    .S(net424),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _11981_ (.A0(net1350),
    .A1(net680),
    .S(net424),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _11982_ (.A0(net1980),
    .A1(net677),
    .S(net424),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(net2472),
    .A1(net676),
    .S(net424),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(net1688),
    .A1(net673),
    .S(net424),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(net2126),
    .A1(net671),
    .S(net424),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _11986_ (.A0(net2752),
    .A1(net668),
    .S(net424),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _11987_ (.A0(net1194),
    .A1(\dpath.RF.wdata[25] ),
    .S(net424),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(net2080),
    .A1(net665),
    .S(net424),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(net1458),
    .A1(net662),
    .S(net424),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _11990_ (.A0(net1266),
    .A1(net661),
    .S(net424),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(net1182),
    .A1(net658),
    .S(net424),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(net3132),
    .A1(net657),
    .S(net424),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(net1264),
    .A1(net655),
    .S(net424),
    .X(_01024_));
 sky130_fd_sc_hd__nand4_1 _11994_ (.A(\ctrl.inst_W[26] ),
    .B(\ctrl.inst_W[27] ),
    .C(\ctrl.inst_W[28] ),
    .D(\ctrl.inst_W[30] ),
    .Y(_05855_));
 sky130_fd_sc_hd__or2_1 _11995_ (.A(\ctrl.inst_W[25] ),
    .B(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__or4b_1 _11996_ (.A(\ctrl.inst_W[31] ),
    .B(\ctrl.inst_W[24] ),
    .C(_02084_),
    .D_N(\ctrl.inst_W[29] ),
    .X(_05857_));
 sky130_fd_sc_hd__or4_4 _11997_ (.A(_01773_),
    .B(_01814_),
    .C(_05856_),
    .D(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__or2_2 _11998_ (.A(\ctrl.inst_W[20] ),
    .B(net471),
    .X(_05859_));
 sky130_fd_sc_hd__or4b_4 _11999_ (.A(\ctrl.inst_W[21] ),
    .B(_05859_),
    .C(\ctrl.inst_W[23] ),
    .D_N(\ctrl.inst_W[22] ),
    .X(_05860_));
 sky130_fd_sc_hd__mux2_1 _12000_ (.A0(net3214),
    .A1(net3571),
    .S(net462),
    .X(_05861_));
 sky130_fd_sc_hd__and2_1 _12001_ (.A(net878),
    .B(net3572),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(net3257),
    .A1(net3560),
    .S(net462),
    .X(_05862_));
 sky130_fd_sc_hd__and2_1 _12003_ (.A(net878),
    .B(net3561),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(net3443),
    .A1(net3603),
    .S(net462),
    .X(_05863_));
 sky130_fd_sc_hd__and2_1 _12005_ (.A(net875),
    .B(net3604),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(net3481),
    .A1(net3563),
    .S(net462),
    .X(_05864_));
 sky130_fd_sc_hd__and2_1 _12007_ (.A(net878),
    .B(net3564),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _12008_ (.A0(net3523),
    .A1(net3566),
    .S(net461),
    .X(_05865_));
 sky130_fd_sc_hd__and2_1 _12009_ (.A(net878),
    .B(_05865_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _12010_ (.A0(net3516),
    .A1(net3557),
    .S(net461),
    .X(_05866_));
 sky130_fd_sc_hd__and2_1 _12011_ (.A(net878),
    .B(_05866_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(net3548),
    .A1(net3562),
    .S(net461),
    .X(_05867_));
 sky130_fd_sc_hd__and2_1 _12013_ (.A(net878),
    .B(_05867_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(net3529),
    .A1(net3554),
    .S(net461),
    .X(_05868_));
 sky130_fd_sc_hd__and2_1 _12015_ (.A(net877),
    .B(_05868_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(net3497),
    .A1(net3553),
    .S(net461),
    .X(_05869_));
 sky130_fd_sc_hd__and2_1 _12017_ (.A(net877),
    .B(_05869_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _12018_ (.A0(net3502),
    .A1(net3581),
    .S(net461),
    .X(_05870_));
 sky130_fd_sc_hd__and2_1 _12019_ (.A(net877),
    .B(_05870_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _12020_ (.A0(net3512),
    .A1(net3577),
    .S(net462),
    .X(_05871_));
 sky130_fd_sc_hd__and2_1 _12021_ (.A(net877),
    .B(net3578),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(\dpath.csrw_out0.d[11] ),
    .A1(net3551),
    .S(net461),
    .X(_05872_));
 sky130_fd_sc_hd__and2_1 _12023_ (.A(net877),
    .B(net3552),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _12024_ (.A0(\dpath.csrw_out0.d[12] ),
    .A1(net3567),
    .S(net461),
    .X(_05873_));
 sky130_fd_sc_hd__and2_1 _12025_ (.A(net877),
    .B(net3568),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _12026_ (.A0(net3433),
    .A1(net3619),
    .S(net462),
    .X(_05874_));
 sky130_fd_sc_hd__and2_1 _12027_ (.A(net878),
    .B(net3620),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _12028_ (.A0(net3457),
    .A1(net3613),
    .S(net462),
    .X(_05875_));
 sky130_fd_sc_hd__and2_1 _12029_ (.A(net878),
    .B(net3614),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _12030_ (.A0(net3404),
    .A1(net3569),
    .S(net462),
    .X(_05876_));
 sky130_fd_sc_hd__and2_1 _12031_ (.A(net875),
    .B(net3570),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(net3366),
    .A1(net3445),
    .S(net462),
    .X(_05877_));
 sky130_fd_sc_hd__and2_1 _12033_ (.A(net875),
    .B(net3446),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _12034_ (.A0(net3334),
    .A1(net3573),
    .S(net462),
    .X(_05878_));
 sky130_fd_sc_hd__and2_1 _12035_ (.A(net875),
    .B(net3574),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(net3247),
    .A1(net3305),
    .S(net462),
    .X(_05879_));
 sky130_fd_sc_hd__and2_1 _12037_ (.A(net875),
    .B(net3306),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _12038_ (.A0(net3488),
    .A1(net3607),
    .S(net461),
    .X(_05880_));
 sky130_fd_sc_hd__and2_1 _12039_ (.A(net877),
    .B(_05880_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _12040_ (.A0(net3486),
    .A1(net3585),
    .S(net461),
    .X(_05881_));
 sky130_fd_sc_hd__and2_1 _12041_ (.A(net877),
    .B(_05881_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _12042_ (.A0(net3500),
    .A1(net3595),
    .S(net461),
    .X(_05882_));
 sky130_fd_sc_hd__and2_1 _12043_ (.A(net877),
    .B(_05882_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _12044_ (.A0(net3448),
    .A1(net3600),
    .S(net461),
    .X(_05883_));
 sky130_fd_sc_hd__and2_1 _12045_ (.A(net877),
    .B(_05883_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _12046_ (.A0(net3255),
    .A1(net3593),
    .S(net461),
    .X(_05884_));
 sky130_fd_sc_hd__and2_1 _12047_ (.A(net877),
    .B(_05884_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(net3217),
    .A1(net3599),
    .S(net461),
    .X(_05885_));
 sky130_fd_sc_hd__and2_1 _12049_ (.A(net878),
    .B(_05885_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(net3450),
    .A1(net3615),
    .S(net462),
    .X(_05886_));
 sky130_fd_sc_hd__and2_1 _12051_ (.A(net877),
    .B(net3616),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(net3430),
    .A1(net3611),
    .S(net462),
    .X(_05887_));
 sky130_fd_sc_hd__and2_1 _12053_ (.A(net877),
    .B(net3612),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _12054_ (.A0(net3380),
    .A1(net3594),
    .S(net461),
    .X(_05888_));
 sky130_fd_sc_hd__and2_1 _12055_ (.A(net877),
    .B(_05888_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _12056_ (.A0(net3459),
    .A1(net3617),
    .S(_05860_),
    .X(_05889_));
 sky130_fd_sc_hd__and2_1 _12057_ (.A(net877),
    .B(net3618),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _12058_ (.A0(net3437),
    .A1(net3608),
    .S(net461),
    .X(_05890_));
 sky130_fd_sc_hd__and2_1 _12059_ (.A(net877),
    .B(_05890_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _12060_ (.A0(net3505),
    .A1(net3596),
    .S(net462),
    .X(_05891_));
 sky130_fd_sc_hd__and2_1 _12061_ (.A(net878),
    .B(net3597),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(net3289),
    .A1(net3591),
    .S(net462),
    .X(_05892_));
 sky130_fd_sc_hd__and2_1 _12063_ (.A(net878),
    .B(net3592),
    .X(_01056_));
 sky130_fd_sc_hd__or3b_2 _12064_ (.A(\ctrl.inst_W[23] ),
    .B(\ctrl.inst_W[22] ),
    .C_N(\ctrl.inst_W[21] ),
    .X(_05893_));
 sky130_fd_sc_hd__nor3_1 _12065_ (.A(net489),
    .B(net470),
    .C(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__or4_1 _12066_ (.A(net3214),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05895_));
 sky130_fd_sc_hd__o211a_1 _12067_ (.A1(net3382),
    .A2(net465),
    .B1(_05895_),
    .C1(net870),
    .X(_01057_));
 sky130_fd_sc_hd__or4_1 _12068_ (.A(net3257),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05896_));
 sky130_fd_sc_hd__o211a_1 _12069_ (.A1(net3406),
    .A2(net465),
    .B1(_05896_),
    .C1(net869),
    .X(_01058_));
 sky130_fd_sc_hd__or4_1 _12070_ (.A(\dpath.csrw_out0.d[2] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05897_));
 sky130_fd_sc_hd__o211a_1 _12071_ (.A1(net3376),
    .A2(net465),
    .B1(_05897_),
    .C1(net870),
    .X(_01059_));
 sky130_fd_sc_hd__or4_1 _12072_ (.A(\dpath.csrw_out0.d[3] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05898_));
 sky130_fd_sc_hd__o211a_1 _12073_ (.A1(net3408),
    .A2(net465),
    .B1(_05898_),
    .C1(net870),
    .X(_01060_));
 sky130_fd_sc_hd__or4_1 _12074_ (.A(\dpath.csrw_out0.d[4] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05899_));
 sky130_fd_sc_hd__o211a_1 _12075_ (.A1(net3347),
    .A2(net465),
    .B1(_05899_),
    .C1(net870),
    .X(_01061_));
 sky130_fd_sc_hd__or4_1 _12076_ (.A(\dpath.csrw_out0.d[5] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05900_));
 sky130_fd_sc_hd__o211a_1 _12077_ (.A1(net3390),
    .A2(net465),
    .B1(_05900_),
    .C1(net870),
    .X(_01062_));
 sky130_fd_sc_hd__or4_1 _12078_ (.A(\dpath.csrw_out0.d[6] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05901_));
 sky130_fd_sc_hd__o211a_1 _12079_ (.A1(net3328),
    .A2(net465),
    .B1(_05901_),
    .C1(net869),
    .X(_01063_));
 sky130_fd_sc_hd__or4_1 _12080_ (.A(\dpath.csrw_out0.d[7] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05902_));
 sky130_fd_sc_hd__o211a_1 _12081_ (.A1(net3343),
    .A2(net465),
    .B1(_05902_),
    .C1(net873),
    .X(_01064_));
 sky130_fd_sc_hd__or4_1 _12082_ (.A(\dpath.csrw_out0.d[8] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05903_));
 sky130_fd_sc_hd__o211a_1 _12083_ (.A1(net3330),
    .A2(net465),
    .B1(_05903_),
    .C1(net873),
    .X(_01065_));
 sky130_fd_sc_hd__or4_1 _12084_ (.A(\dpath.csrw_out0.d[9] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05904_));
 sky130_fd_sc_hd__o211a_1 _12085_ (.A1(net3364),
    .A2(net465),
    .B1(_05904_),
    .C1(net873),
    .X(_01066_));
 sky130_fd_sc_hd__or4_1 _12086_ (.A(\dpath.csrw_out0.d[10] ),
    .B(net490),
    .C(_05858_),
    .D(net487),
    .X(_05905_));
 sky130_fd_sc_hd__o211a_1 _12087_ (.A1(net3352),
    .A2(net466),
    .B1(_05905_),
    .C1(net873),
    .X(_01067_));
 sky130_fd_sc_hd__or4_1 _12088_ (.A(\dpath.csrw_out0.d[11] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05906_));
 sky130_fd_sc_hd__o211a_1 _12089_ (.A1(net3319),
    .A2(net465),
    .B1(_05906_),
    .C1(net873),
    .X(_01068_));
 sky130_fd_sc_hd__or4_1 _12090_ (.A(\dpath.csrw_out0.d[12] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05907_));
 sky130_fd_sc_hd__o211a_1 _12091_ (.A1(net3317),
    .A2(net465),
    .B1(_05907_),
    .C1(net873),
    .X(_01069_));
 sky130_fd_sc_hd__or4_1 _12092_ (.A(\dpath.csrw_out0.d[13] ),
    .B(net489),
    .C(net470),
    .D(net487),
    .X(_05908_));
 sky130_fd_sc_hd__o211a_1 _12093_ (.A1(net3315),
    .A2(net465),
    .B1(_05908_),
    .C1(net873),
    .X(_01070_));
 sky130_fd_sc_hd__or4_1 _12094_ (.A(\dpath.csrw_out0.d[14] ),
    .B(net489),
    .C(net470),
    .D(_05893_),
    .X(_05909_));
 sky130_fd_sc_hd__o211a_1 _12095_ (.A1(net3313),
    .A2(net465),
    .B1(_05909_),
    .C1(net873),
    .X(_01071_));
 sky130_fd_sc_hd__or4_1 _12096_ (.A(\dpath.csrw_out0.d[15] ),
    .B(net489),
    .C(net470),
    .D(net488),
    .X(_05910_));
 sky130_fd_sc_hd__o211a_1 _12097_ (.A1(net3293),
    .A2(net465),
    .B1(_05910_),
    .C1(net873),
    .X(_01072_));
 sky130_fd_sc_hd__or4_1 _12098_ (.A(\dpath.csrw_out0.d[16] ),
    .B(_01791_),
    .C(net471),
    .D(net488),
    .X(_05911_));
 sky130_fd_sc_hd__o211a_1 _12099_ (.A1(net3299),
    .A2(net465),
    .B1(_05911_),
    .C1(net874),
    .X(_01073_));
 sky130_fd_sc_hd__or4_1 _12100_ (.A(\dpath.csrw_out0.d[17] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05912_));
 sky130_fd_sc_hd__o211a_1 _12101_ (.A1(net3332),
    .A2(net466),
    .B1(_05912_),
    .C1(net875),
    .X(_01074_));
 sky130_fd_sc_hd__or4_1 _12102_ (.A(net3247),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05913_));
 sky130_fd_sc_hd__o211a_1 _12103_ (.A1(net3303),
    .A2(net466),
    .B1(_05913_),
    .C1(net875),
    .X(_01075_));
 sky130_fd_sc_hd__or4_1 _12104_ (.A(\dpath.csrw_out0.d[19] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05914_));
 sky130_fd_sc_hd__o211a_1 _12105_ (.A1(net3321),
    .A2(net466),
    .B1(_05914_),
    .C1(net875),
    .X(_01076_));
 sky130_fd_sc_hd__or4_1 _12106_ (.A(\dpath.csrw_out0.d[20] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05915_));
 sky130_fd_sc_hd__o211a_1 _12107_ (.A1(net3370),
    .A2(net466),
    .B1(_05915_),
    .C1(net875),
    .X(_01077_));
 sky130_fd_sc_hd__or4_1 _12108_ (.A(\dpath.csrw_out0.d[21] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05916_));
 sky130_fd_sc_hd__o211a_1 _12109_ (.A1(net3350),
    .A2(net466),
    .B1(_05916_),
    .C1(net875),
    .X(_01078_));
 sky130_fd_sc_hd__or4_1 _12110_ (.A(\dpath.csrw_out0.d[22] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05917_));
 sky130_fd_sc_hd__o211a_1 _12111_ (.A1(net3360),
    .A2(_05894_),
    .B1(_05917_),
    .C1(net875),
    .X(_01079_));
 sky130_fd_sc_hd__or4_1 _12112_ (.A(net3255),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05918_));
 sky130_fd_sc_hd__o211a_1 _12113_ (.A1(net3362),
    .A2(net466),
    .B1(_05918_),
    .C1(net875),
    .X(_01080_));
 sky130_fd_sc_hd__or4_1 _12114_ (.A(net3217),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05919_));
 sky130_fd_sc_hd__o211a_1 _12115_ (.A1(net3354),
    .A2(net466),
    .B1(_05919_),
    .C1(net875),
    .X(_01081_));
 sky130_fd_sc_hd__or4_1 _12116_ (.A(\dpath.csrw_out0.d[25] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05920_));
 sky130_fd_sc_hd__o211a_1 _12117_ (.A1(net3356),
    .A2(net466),
    .B1(_05920_),
    .C1(net875),
    .X(_01082_));
 sky130_fd_sc_hd__or4_1 _12118_ (.A(\dpath.csrw_out0.d[26] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05921_));
 sky130_fd_sc_hd__o211a_1 _12119_ (.A1(net3388),
    .A2(net466),
    .B1(_05921_),
    .C1(net876),
    .X(_01083_));
 sky130_fd_sc_hd__or4_1 _12120_ (.A(net3380),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05922_));
 sky130_fd_sc_hd__o211a_1 _12121_ (.A1(net3386),
    .A2(net466),
    .B1(_05922_),
    .C1(net875),
    .X(_01084_));
 sky130_fd_sc_hd__or4_1 _12122_ (.A(\dpath.csrw_out0.d[28] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05923_));
 sky130_fd_sc_hd__o211a_1 _12123_ (.A1(net3384),
    .A2(net466),
    .B1(_05923_),
    .C1(net878),
    .X(_01085_));
 sky130_fd_sc_hd__or4_1 _12124_ (.A(\dpath.csrw_out0.d[29] ),
    .B(net490),
    .C(net471),
    .D(_05893_),
    .X(_05924_));
 sky130_fd_sc_hd__o211a_1 _12125_ (.A1(net3413),
    .A2(net466),
    .B1(_05924_),
    .C1(net878),
    .X(_01086_));
 sky130_fd_sc_hd__or4_1 _12126_ (.A(\dpath.csrw_out0.d[30] ),
    .B(net490),
    .C(net471),
    .D(net488),
    .X(_05925_));
 sky130_fd_sc_hd__o211a_1 _12127_ (.A1(net3378),
    .A2(net466),
    .B1(_05925_),
    .C1(net878),
    .X(_01087_));
 sky130_fd_sc_hd__or4_1 _12128_ (.A(net3289),
    .B(_01791_),
    .C(_05858_),
    .D(net488),
    .X(_05926_));
 sky130_fd_sc_hd__o211a_1 _12129_ (.A1(net3418),
    .A2(net466),
    .B1(_05926_),
    .C1(net878),
    .X(_01088_));
 sky130_fd_sc_hd__nor2_1 _12130_ (.A(_05859_),
    .B(net487),
    .Y(_05927_));
 sky130_fd_sc_hd__or2_1 _12131_ (.A(_05859_),
    .B(net487),
    .X(_05928_));
 sky130_fd_sc_hd__or2_1 _12132_ (.A(net260),
    .B(net460),
    .X(_05929_));
 sky130_fd_sc_hd__o211a_1 _12133_ (.A1(net3214),
    .A2(net458),
    .B1(_05929_),
    .C1(net869),
    .X(_01089_));
 sky130_fd_sc_hd__or2_1 _12134_ (.A(net271),
    .B(net460),
    .X(_05930_));
 sky130_fd_sc_hd__o211a_1 _12135_ (.A1(net3257),
    .A2(net458),
    .B1(_05930_),
    .C1(net869),
    .X(_01090_));
 sky130_fd_sc_hd__or2_1 _12136_ (.A(net282),
    .B(net460),
    .X(_05931_));
 sky130_fd_sc_hd__o211a_1 _12137_ (.A1(net3443),
    .A2(net458),
    .B1(_05931_),
    .C1(net866),
    .X(_01091_));
 sky130_fd_sc_hd__or2_1 _12138_ (.A(net285),
    .B(net460),
    .X(_05932_));
 sky130_fd_sc_hd__o211a_1 _12139_ (.A1(net3481),
    .A2(net458),
    .B1(_05932_),
    .C1(net866),
    .X(_01092_));
 sky130_fd_sc_hd__or2_1 _12140_ (.A(net286),
    .B(net459),
    .X(_05933_));
 sky130_fd_sc_hd__o211a_1 _12141_ (.A1(net3523),
    .A2(net457),
    .B1(_05933_),
    .C1(net872),
    .X(_01093_));
 sky130_fd_sc_hd__or2_1 _12142_ (.A(net287),
    .B(net459),
    .X(_05934_));
 sky130_fd_sc_hd__o211a_1 _12143_ (.A1(net3516),
    .A2(net457),
    .B1(_05934_),
    .C1(net872),
    .X(_01094_));
 sky130_fd_sc_hd__or2_1 _12144_ (.A(net288),
    .B(net459),
    .X(_05935_));
 sky130_fd_sc_hd__o211a_1 _12145_ (.A1(net3548),
    .A2(net457),
    .B1(_05935_),
    .C1(net872),
    .X(_01095_));
 sky130_fd_sc_hd__or2_1 _12146_ (.A(net289),
    .B(net459),
    .X(_05936_));
 sky130_fd_sc_hd__o211a_1 _12147_ (.A1(net3529),
    .A2(net457),
    .B1(_05936_),
    .C1(net872),
    .X(_01096_));
 sky130_fd_sc_hd__or2_1 _12148_ (.A(net290),
    .B(net459),
    .X(_05937_));
 sky130_fd_sc_hd__o211a_1 _12149_ (.A1(net3497),
    .A2(net457),
    .B1(_05937_),
    .C1(net866),
    .X(_01097_));
 sky130_fd_sc_hd__or2_1 _12150_ (.A(net291),
    .B(net459),
    .X(_05938_));
 sky130_fd_sc_hd__o211a_1 _12151_ (.A1(net3502),
    .A2(net457),
    .B1(_05938_),
    .C1(net872),
    .X(_01098_));
 sky130_fd_sc_hd__or2_1 _12152_ (.A(net261),
    .B(net459),
    .X(_05939_));
 sky130_fd_sc_hd__o211a_1 _12153_ (.A1(net3512),
    .A2(net457),
    .B1(_05939_),
    .C1(net872),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _12154_ (.A(net3520),
    .B(net459),
    .X(_05940_));
 sky130_fd_sc_hd__o211a_1 _12155_ (.A1(\dpath.csrw_out0.d[11] ),
    .A2(net457),
    .B1(_05940_),
    .C1(net872),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _12156_ (.A(net3532),
    .B(net459),
    .X(_05941_));
 sky130_fd_sc_hd__o211a_1 _12157_ (.A1(\dpath.csrw_out0.d[12] ),
    .A2(net457),
    .B1(_05941_),
    .C1(net872),
    .X(_01101_));
 sky130_fd_sc_hd__or2_1 _12158_ (.A(net264),
    .B(net460),
    .X(_05942_));
 sky130_fd_sc_hd__o211a_1 _12159_ (.A1(net3433),
    .A2(net458),
    .B1(_05942_),
    .C1(net867),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _12160_ (.A(net265),
    .B(net459),
    .X(_05943_));
 sky130_fd_sc_hd__o211a_1 _12161_ (.A1(net3457),
    .A2(net457),
    .B1(_05943_),
    .C1(net872),
    .X(_01103_));
 sky130_fd_sc_hd__or2_1 _12162_ (.A(net266),
    .B(net459),
    .X(_05944_));
 sky130_fd_sc_hd__o211a_1 _12163_ (.A1(net3404),
    .A2(net457),
    .B1(_05944_),
    .C1(net872),
    .X(_01104_));
 sky130_fd_sc_hd__or2_1 _12164_ (.A(net267),
    .B(net459),
    .X(_05945_));
 sky130_fd_sc_hd__o211a_1 _12165_ (.A1(net3366),
    .A2(net457),
    .B1(_05945_),
    .C1(net866),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _12166_ (.A(net268),
    .B(net459),
    .X(_05946_));
 sky130_fd_sc_hd__o211a_1 _12167_ (.A1(net3334),
    .A2(net457),
    .B1(_05946_),
    .C1(net866),
    .X(_01106_));
 sky130_fd_sc_hd__or2_1 _12168_ (.A(net269),
    .B(net459),
    .X(_05947_));
 sky130_fd_sc_hd__o211a_1 _12169_ (.A1(net3247),
    .A2(net457),
    .B1(_05947_),
    .C1(net866),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _12170_ (.A(net270),
    .B(net459),
    .X(_05948_));
 sky130_fd_sc_hd__o211a_1 _12171_ (.A1(net3488),
    .A2(net457),
    .B1(_05948_),
    .C1(net866),
    .X(_01108_));
 sky130_fd_sc_hd__or2_1 _12172_ (.A(net272),
    .B(net459),
    .X(_05949_));
 sky130_fd_sc_hd__o211a_1 _12173_ (.A1(net3486),
    .A2(net457),
    .B1(_05949_),
    .C1(net866),
    .X(_01109_));
 sky130_fd_sc_hd__or2_1 _12174_ (.A(net273),
    .B(net460),
    .X(_05950_));
 sky130_fd_sc_hd__o211a_1 _12175_ (.A1(net3500),
    .A2(net458),
    .B1(_05950_),
    .C1(net866),
    .X(_01110_));
 sky130_fd_sc_hd__or2_1 _12176_ (.A(net274),
    .B(net460),
    .X(_05951_));
 sky130_fd_sc_hd__o211a_1 _12177_ (.A1(net3448),
    .A2(net458),
    .B1(_05951_),
    .C1(net867),
    .X(_01111_));
 sky130_fd_sc_hd__or2_1 _12178_ (.A(net275),
    .B(_05927_),
    .X(_05952_));
 sky130_fd_sc_hd__o211a_1 _12179_ (.A1(net3255),
    .A2(_05928_),
    .B1(_05952_),
    .C1(net867),
    .X(_01112_));
 sky130_fd_sc_hd__or2_1 _12180_ (.A(net276),
    .B(net460),
    .X(_05953_));
 sky130_fd_sc_hd__o211a_1 _12181_ (.A1(net3217),
    .A2(net458),
    .B1(_05953_),
    .C1(net867),
    .X(_01113_));
 sky130_fd_sc_hd__or2_1 _12182_ (.A(net277),
    .B(net460),
    .X(_05954_));
 sky130_fd_sc_hd__o211a_1 _12183_ (.A1(net3450),
    .A2(net458),
    .B1(_05954_),
    .C1(net867),
    .X(_01114_));
 sky130_fd_sc_hd__or2_1 _12184_ (.A(net278),
    .B(net460),
    .X(_05955_));
 sky130_fd_sc_hd__o211a_1 _12185_ (.A1(net3430),
    .A2(net458),
    .B1(_05955_),
    .C1(net869),
    .X(_01115_));
 sky130_fd_sc_hd__or2_1 _12186_ (.A(net279),
    .B(net460),
    .X(_05956_));
 sky130_fd_sc_hd__o211a_1 _12187_ (.A1(net3380),
    .A2(net458),
    .B1(_05956_),
    .C1(net869),
    .X(_01116_));
 sky130_fd_sc_hd__or2_1 _12188_ (.A(net280),
    .B(net460),
    .X(_05957_));
 sky130_fd_sc_hd__o211a_1 _12189_ (.A1(net3459),
    .A2(net458),
    .B1(_05957_),
    .C1(net869),
    .X(_01117_));
 sky130_fd_sc_hd__or2_1 _12190_ (.A(net281),
    .B(net460),
    .X(_05958_));
 sky130_fd_sc_hd__o211a_1 _12191_ (.A1(net3437),
    .A2(net458),
    .B1(_05958_),
    .C1(net869),
    .X(_01118_));
 sky130_fd_sc_hd__or2_1 _12192_ (.A(net283),
    .B(net460),
    .X(_05959_));
 sky130_fd_sc_hd__o211a_1 _12193_ (.A1(net3505),
    .A2(net458),
    .B1(_05959_),
    .C1(net869),
    .X(_01119_));
 sky130_fd_sc_hd__or2_1 _12194_ (.A(net284),
    .B(net460),
    .X(_05960_));
 sky130_fd_sc_hd__o211a_1 _12195_ (.A1(net3289),
    .A2(net458),
    .B1(_05960_),
    .C1(net869),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _12196_ (.A0(\dpath.RF.R[4][0] ),
    .A1(\dpath.RF.R[5][0] ),
    .A2(\dpath.RF.R[6][0] ),
    .A3(\dpath.RF.R[7][0] ),
    .S0(net563),
    .S1(net546),
    .X(_05961_));
 sky130_fd_sc_hd__mux2_1 _12197_ (.A0(\dpath.RF.R[0][0] ),
    .A1(\dpath.RF.R[1][0] ),
    .S(net563),
    .X(_05962_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(\dpath.RF.R[2][0] ),
    .A1(\dpath.RF.R[3][0] ),
    .S(net563),
    .X(_05963_));
 sky130_fd_sc_hd__a21o_1 _12199_ (.A1(net546),
    .A2(_05963_),
    .B1(net531),
    .X(_05964_));
 sky130_fd_sc_hd__a21o_1 _12200_ (.A1(_01770_),
    .A2(_05962_),
    .B1(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__o211a_1 _12201_ (.A1(net511),
    .A2(_05961_),
    .B1(_05965_),
    .C1(net506),
    .X(_05966_));
 sky130_fd_sc_hd__mux4_1 _12202_ (.A0(\dpath.RF.R[8][0] ),
    .A1(\dpath.RF.R[9][0] ),
    .A2(\dpath.RF.R[10][0] ),
    .A3(\dpath.RF.R[11][0] ),
    .S0(net562),
    .S1(net543),
    .X(_05967_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(\dpath.RF.R[14][0] ),
    .A1(\dpath.RF.R[15][0] ),
    .S(net562),
    .X(_05968_));
 sky130_fd_sc_hd__mux2_1 _12204_ (.A0(\dpath.RF.R[12][0] ),
    .A1(\dpath.RF.R[13][0] ),
    .S(net562),
    .X(_05969_));
 sky130_fd_sc_hd__a21o_1 _12205_ (.A1(_01770_),
    .A2(_05969_),
    .B1(net511),
    .X(_05970_));
 sky130_fd_sc_hd__a21o_1 _12206_ (.A1(net543),
    .A2(_05968_),
    .B1(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__o211a_1 _12207_ (.A1(net531),
    .A2(_05967_),
    .B1(_05971_),
    .C1(net523),
    .X(_05972_));
 sky130_fd_sc_hd__or3_1 _12208_ (.A(net518),
    .B(_05966_),
    .C(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__mux4_1 _12209_ (.A0(\dpath.RF.R[16][0] ),
    .A1(\dpath.RF.R[17][0] ),
    .A2(\dpath.RF.R[18][0] ),
    .A3(\dpath.RF.R[19][0] ),
    .S0(net563),
    .S1(net546),
    .X(_05974_));
 sky130_fd_sc_hd__nor2_1 _12210_ (.A(net531),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__mux4_1 _12211_ (.A0(\dpath.RF.R[20][0] ),
    .A1(\dpath.RF.R[21][0] ),
    .A2(\dpath.RF.R[22][0] ),
    .A3(\dpath.RF.R[23][0] ),
    .S0(net563),
    .S1(net546),
    .X(_05976_));
 sky130_fd_sc_hd__nor2_1 _12212_ (.A(net511),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__mux4_1 _12213_ (.A0(\dpath.RF.R[28][0] ),
    .A1(\dpath.RF.R[29][0] ),
    .A2(\dpath.RF.R[30][0] ),
    .A3(\dpath.RF.R[31][0] ),
    .S0(net562),
    .S1(net543),
    .X(_05978_));
 sky130_fd_sc_hd__nor2_1 _12214_ (.A(net511),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__mux4_1 _12215_ (.A0(\dpath.RF.R[24][0] ),
    .A1(\dpath.RF.R[25][0] ),
    .A2(\dpath.RF.R[26][0] ),
    .A3(\dpath.RF.R[27][0] ),
    .S0(net563),
    .S1(net543),
    .X(_05980_));
 sky130_fd_sc_hd__o21ai_1 _12216_ (.A1(net531),
    .A2(_05980_),
    .B1(net523),
    .Y(_05981_));
 sky130_fd_sc_hd__o32a_1 _12217_ (.A1(net523),
    .A2(_05975_),
    .A3(_05977_),
    .B1(_05979_),
    .B2(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__nand2_1 _12218_ (.A(net518),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__and4bb_1 _12219_ (.A_N(net482),
    .B_N(net372),
    .C(_05973_),
    .D(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(net3652),
    .A1(_01842_),
    .S(net484),
    .X(_05985_));
 sky130_fd_sc_hd__nand2_1 _12221_ (.A(_01951_),
    .B(net467),
    .Y(_05986_));
 sky130_fd_sc_hd__o21ai_4 _12222_ (.A1(net467),
    .A2(_05985_),
    .B1(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__mux2_4 _12224_ (.A0(net3605),
    .A1(net1),
    .S(net480),
    .X(_05989_));
 sky130_fd_sc_hd__a221o_1 _12225_ (.A1(net392),
    .A2(_05988_),
    .B1(_05989_),
    .B2(net368),
    .C1(_05984_),
    .X(_05990_));
 sky130_fd_sc_hd__a21oi_4 _12226_ (.A1(net719),
    .A2(net370),
    .B1(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__nor2_2 _12227_ (.A(net882),
    .B(_05991_),
    .Y(_01121_));
 sky130_fd_sc_hd__mux4_1 _12228_ (.A0(\dpath.RF.R[0][1] ),
    .A1(\dpath.RF.R[1][1] ),
    .A2(\dpath.RF.R[2][1] ),
    .A3(\dpath.RF.R[3][1] ),
    .S0(net562),
    .S1(net543),
    .X(_05992_));
 sky130_fd_sc_hd__nor2_1 _12229_ (.A(net531),
    .B(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__mux2_1 _12230_ (.A0(\dpath.RF.R[6][1] ),
    .A1(\dpath.RF.R[7][1] ),
    .S(net562),
    .X(_05994_));
 sky130_fd_sc_hd__nand2_1 _12231_ (.A(net543),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(\dpath.RF.R[4][1] ),
    .A1(\dpath.RF.R[5][1] ),
    .S(net562),
    .X(_05996_));
 sky130_fd_sc_hd__nand2_1 _12233_ (.A(_01770_),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__a311o_1 _12234_ (.A1(net531),
    .A2(_05995_),
    .A3(_05997_),
    .B1(net523),
    .C1(_05993_),
    .X(_05998_));
 sky130_fd_sc_hd__mux4_1 _12235_ (.A0(\dpath.RF.R[12][1] ),
    .A1(\dpath.RF.R[13][1] ),
    .A2(\dpath.RF.R[14][1] ),
    .A3(\dpath.RF.R[15][1] ),
    .S0(net562),
    .S1(net543),
    .X(_05999_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(\dpath.RF.R[8][1] ),
    .A1(\dpath.RF.R[9][1] ),
    .S(net562),
    .X(_06000_));
 sky130_fd_sc_hd__mux2_1 _12237_ (.A0(\dpath.RF.R[10][1] ),
    .A1(\dpath.RF.R[11][1] ),
    .S(net562),
    .X(_06001_));
 sky130_fd_sc_hd__a21o_1 _12238_ (.A1(net543),
    .A2(_06001_),
    .B1(net531),
    .X(_06002_));
 sky130_fd_sc_hd__a21o_1 _12239_ (.A1(_01770_),
    .A2(_06000_),
    .B1(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__o211a_1 _12240_ (.A1(net511),
    .A2(_05999_),
    .B1(_06003_),
    .C1(net523),
    .X(_06004_));
 sky130_fd_sc_hd__nor2_1 _12241_ (.A(net518),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__mux4_1 _12242_ (.A0(\dpath.RF.R[16][1] ),
    .A1(\dpath.RF.R[17][1] ),
    .A2(\dpath.RF.R[18][1] ),
    .A3(\dpath.RF.R[19][1] ),
    .S0(net562),
    .S1(net543),
    .X(_06006_));
 sky130_fd_sc_hd__nor2_1 _12243_ (.A(net531),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__mux4_1 _12244_ (.A0(\dpath.RF.R[20][1] ),
    .A1(\dpath.RF.R[21][1] ),
    .A2(\dpath.RF.R[22][1] ),
    .A3(\dpath.RF.R[23][1] ),
    .S0(net565),
    .S1(net544),
    .X(_06008_));
 sky130_fd_sc_hd__nor2_1 _12245_ (.A(net511),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__mux4_1 _12246_ (.A0(\dpath.RF.R[28][1] ),
    .A1(\dpath.RF.R[29][1] ),
    .A2(\dpath.RF.R[30][1] ),
    .A3(\dpath.RF.R[31][1] ),
    .S0(net562),
    .S1(net543),
    .X(_06010_));
 sky130_fd_sc_hd__nor2_1 _12247_ (.A(net511),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__mux4_1 _12248_ (.A0(\dpath.RF.R[24][1] ),
    .A1(\dpath.RF.R[25][1] ),
    .A2(\dpath.RF.R[26][1] ),
    .A3(\dpath.RF.R[27][1] ),
    .S0(net562),
    .S1(net543),
    .X(_06012_));
 sky130_fd_sc_hd__o21ai_1 _12249_ (.A1(net531),
    .A2(_06012_),
    .B1(net523),
    .Y(_06013_));
 sky130_fd_sc_hd__o32a_1 _12250_ (.A1(net523),
    .A2(_06007_),
    .A3(_06009_),
    .B1(_06011_),
    .B2(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__a22o_1 _12251_ (.A1(_05998_),
    .A2(_06005_),
    .B1(_06014_),
    .B2(net518),
    .X(_06015_));
 sky130_fd_sc_hd__nor3_1 _12252_ (.A(net482),
    .B(net372),
    .C(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__mux2_2 _12253_ (.A0(net3541),
    .A1(net12),
    .S(net480),
    .X(_06017_));
 sky130_fd_sc_hd__xor2_1 _12254_ (.A(_01842_),
    .B(_01905_),
    .X(_06018_));
 sky130_fd_sc_hd__a22o_1 _12255_ (.A1(net786),
    .A2(net647),
    .B1(net783),
    .B2(net651),
    .X(_06019_));
 sky130_fd_sc_hd__nand2_1 _12256_ (.A(net484),
    .B(_06019_),
    .Y(_06020_));
 sky130_fd_sc_hd__a2bb2o_1 _12257_ (.A1_N(_02108_),
    .A2_N(_06020_),
    .B1(net3682),
    .B2(net485),
    .X(_06021_));
 sky130_fd_sc_hd__mux2_4 _12258_ (.A0(_06018_),
    .A1(_06021_),
    .S(net468),
    .X(_06022_));
 sky130_fd_sc_hd__a22o_1 _12259_ (.A1(net368),
    .A2(_06017_),
    .B1(_06022_),
    .B2(net392),
    .X(_06023_));
 sky130_fd_sc_hd__a211o_2 _12260_ (.A1(net716),
    .A2(net370),
    .B1(_06016_),
    .C1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__and2_1 _12261_ (.A(net862),
    .B(_06024_),
    .X(_01122_));
 sky130_fd_sc_hd__and2_1 _12262_ (.A(net849),
    .B(_02118_),
    .X(_01123_));
 sky130_fd_sc_hd__nor2_1 _12263_ (.A(net883),
    .B(net3273),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _12264_ (.A(net882),
    .B(net3269),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _12265_ (.A(net888),
    .B(_02317_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _12266_ (.A(net882),
    .B(net3412),
    .Y(_01127_));
 sky130_fd_sc_hd__nor2_1 _12267_ (.A(net888),
    .B(net3400),
    .Y(_01128_));
 sky130_fd_sc_hd__nor2_2 _12268_ (.A(net888),
    .B(_02552_),
    .Y(_01129_));
 sky130_fd_sc_hd__nor2_1 _12269_ (.A(net887),
    .B(_02641_),
    .Y(_01130_));
 sky130_fd_sc_hd__nor2_2 _12270_ (.A(net888),
    .B(_02741_),
    .Y(_01131_));
 sky130_fd_sc_hd__nor2_1 _12271_ (.A(net888),
    .B(net3629),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_2 _12272_ (.A(net888),
    .B(_02945_),
    .Y(_01133_));
 sky130_fd_sc_hd__and2_1 _12273_ (.A(net871),
    .B(_03053_),
    .X(_01134_));
 sky130_fd_sc_hd__nor2_2 _12274_ (.A(net888),
    .B(_03167_),
    .Y(_01135_));
 sky130_fd_sc_hd__and2_1 _12275_ (.A(net871),
    .B(_03283_),
    .X(_01136_));
 sky130_fd_sc_hd__nor2_2 _12276_ (.A(net884),
    .B(_03412_),
    .Y(_01137_));
 sky130_fd_sc_hd__and2_1 _12277_ (.A(net871),
    .B(_03544_),
    .X(_01138_));
 sky130_fd_sc_hd__nor2_2 _12278_ (.A(net884),
    .B(_03685_),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_2 _12279_ (.A(net887),
    .B(_03821_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_2 _12280_ (.A(net887),
    .B(_03969_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_2 _12281_ (.A(net887),
    .B(_04114_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_2 _12282_ (.A(net887),
    .B(_04276_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_2 _12283_ (.A(net885),
    .B(_04422_),
    .Y(_01144_));
 sky130_fd_sc_hd__and2_2 _12284_ (.A(net879),
    .B(_04594_),
    .X(_01145_));
 sky130_fd_sc_hd__nor2_2 _12285_ (.A(net885),
    .B(_04760_),
    .Y(_01146_));
 sky130_fd_sc_hd__and2_2 _12286_ (.A(net862),
    .B(_04934_),
    .X(_01147_));
 sky130_fd_sc_hd__nor2_1 _12287_ (.A(net885),
    .B(_05110_),
    .Y(_01148_));
 sky130_fd_sc_hd__and2_1 _12288_ (.A(net879),
    .B(_05293_),
    .X(_01149_));
 sky130_fd_sc_hd__nor2_1 _12289_ (.A(net885),
    .B(_05477_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_2 _12290_ (.A(net886),
    .B(_05663_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _12291_ (.A(net885),
    .B(_05829_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _12292_ (.A(\ctrl.d2c_inst[23] ),
    .B(\ctrl.d2c_inst[22] ),
    .Y(_06025_));
 sky130_fd_sc_hd__nor2_1 _12293_ (.A(\ctrl.d2c_inst[21] ),
    .B(\ctrl.d2c_inst[20] ),
    .Y(_06026_));
 sky130_fd_sc_hd__and3_1 _12294_ (.A(_01749_),
    .B(_06025_),
    .C(_06026_),
    .X(_06027_));
 sky130_fd_sc_hd__a22o_1 _12295_ (.A1(_01752_),
    .A2(\ctrl.c2d_rf_waddr_W[1] ),
    .B1(\ctrl.c2d_rf_waddr_W[4] ),
    .B2(_01749_),
    .X(_06028_));
 sky130_fd_sc_hd__a221o_1 _12296_ (.A1(_01751_),
    .A2(\ctrl.c2d_rf_waddr_W[2] ),
    .B1(_01780_),
    .B2(\ctrl.d2c_inst[24] ),
    .C1(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__a22o_1 _12297_ (.A1(\ctrl.d2c_inst[22] ),
    .A2(_01778_),
    .B1(\ctrl.c2d_rf_waddr_W[3] ),
    .B2(_01750_),
    .X(_06030_));
 sky130_fd_sc_hd__a2111o_1 _12298_ (.A1(\ctrl.d2c_inst[23] ),
    .A2(_01779_),
    .B1(_06029_),
    .C1(_06030_),
    .D1(_01773_),
    .X(_06031_));
 sky130_fd_sc_hd__a22o_1 _12299_ (.A1(\ctrl.d2c_inst[20] ),
    .A2(_01776_),
    .B1(_01777_),
    .B2(\ctrl.d2c_inst[21] ),
    .X(_06032_));
 sky130_fd_sc_hd__a211o_1 _12300_ (.A1(_01753_),
    .A2(\ctrl.c2d_rf_waddr_W[0] ),
    .B1(_02091_),
    .C1(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__or4b_2 _12301_ (.A(_02086_),
    .B(_06031_),
    .C(_06033_),
    .D_N(_01983_),
    .X(_06034_));
 sky130_fd_sc_hd__o22a_1 _12302_ (.A1(_01753_),
    .A2(\ctrl.inst_M[7] ),
    .B1(_01781_),
    .B2(\ctrl.d2c_inst[21] ),
    .X(_06035_));
 sky130_fd_sc_hd__o221a_1 _12303_ (.A1(_01752_),
    .A2(\ctrl.inst_M[8] ),
    .B1(_01782_),
    .B2(\ctrl.d2c_inst[22] ),
    .C1(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__o22a_1 _12304_ (.A1(_01751_),
    .A2(\ctrl.inst_M[9] ),
    .B1(_01784_),
    .B2(\ctrl.d2c_inst[24] ),
    .X(_06037_));
 sky130_fd_sc_hd__o2111a_1 _12305_ (.A1(_01749_),
    .A2(\ctrl.inst_M[11] ),
    .B1(_06036_),
    .C1(_06037_),
    .D1(\ctrl.val_M ),
    .X(_06038_));
 sky130_fd_sc_hd__o2bb2a_1 _12306_ (.A1_N(_01753_),
    .A2_N(\ctrl.inst_M[7] ),
    .B1(\ctrl.inst_M[10] ),
    .B2(_01750_),
    .X(_06039_));
 sky130_fd_sc_hd__o211a_1 _12307_ (.A1(\ctrl.d2c_inst[23] ),
    .A2(_01783_),
    .B1(_02057_),
    .C1(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__and4_1 _12308_ (.A(_01983_),
    .B(_02053_),
    .C(_06038_),
    .D(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__a21oi_1 _12309_ (.A1(_01995_),
    .A2(_02076_),
    .B1(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__and3b_1 _12310_ (.A_N(_06027_),
    .B(_06034_),
    .C(net380),
    .X(_06043_));
 sky130_fd_sc_hd__mux4_1 _12311_ (.A0(\dpath.RF.R[16][0] ),
    .A1(\dpath.RF.R[17][0] ),
    .A2(\dpath.RF.R[18][0] ),
    .A3(\dpath.RF.R[19][0] ),
    .S0(net829),
    .S1(net808),
    .X(_06044_));
 sky130_fd_sc_hd__mux4_1 _12312_ (.A0(\dpath.RF.R[20][0] ),
    .A1(\dpath.RF.R[21][0] ),
    .A2(\dpath.RF.R[22][0] ),
    .A3(\dpath.RF.R[23][0] ),
    .S0(net829),
    .S1(net805),
    .X(_06045_));
 sky130_fd_sc_hd__mux4_1 _12313_ (.A0(\dpath.RF.R[28][0] ),
    .A1(\dpath.RF.R[29][0] ),
    .A2(\dpath.RF.R[30][0] ),
    .A3(\dpath.RF.R[31][0] ),
    .S0(net825),
    .S1(net805),
    .X(_06046_));
 sky130_fd_sc_hd__mux4_1 _12314_ (.A0(\dpath.RF.R[24][0] ),
    .A1(\dpath.RF.R[25][0] ),
    .A2(\dpath.RF.R[26][0] ),
    .A3(\dpath.RF.R[27][0] ),
    .S0(net829),
    .S1(net805),
    .X(_06047_));
 sky130_fd_sc_hd__mux4_1 _12315_ (.A0(_06044_),
    .A1(_06045_),
    .A2(_06047_),
    .A3(_06046_),
    .S0(net797),
    .S1(net794),
    .X(_06048_));
 sky130_fd_sc_hd__inv_2 _12316_ (.A(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__mux4_1 _12317_ (.A0(\dpath.RF.R[12][0] ),
    .A1(\dpath.RF.R[13][0] ),
    .A2(\dpath.RF.R[14][0] ),
    .A3(\dpath.RF.R[15][0] ),
    .S0(net825),
    .S1(net805),
    .X(_06050_));
 sky130_fd_sc_hd__mux4_1 _12318_ (.A0(\dpath.RF.R[8][0] ),
    .A1(\dpath.RF.R[9][0] ),
    .A2(\dpath.RF.R[10][0] ),
    .A3(\dpath.RF.R[11][0] ),
    .S0(net825),
    .S1(net805),
    .X(_06051_));
 sky130_fd_sc_hd__mux4_1 _12319_ (.A0(\dpath.RF.R[0][0] ),
    .A1(\dpath.RF.R[1][0] ),
    .A2(\dpath.RF.R[2][0] ),
    .A3(\dpath.RF.R[3][0] ),
    .S0(net825),
    .S1(net808),
    .X(_06052_));
 sky130_fd_sc_hd__mux4_1 _12320_ (.A0(\dpath.RF.R[4][0] ),
    .A1(\dpath.RF.R[5][0] ),
    .A2(\dpath.RF.R[6][0] ),
    .A3(\dpath.RF.R[7][0] ),
    .S0(net829),
    .S1(net808),
    .X(_06053_));
 sky130_fd_sc_hd__mux4_1 _12321_ (.A0(_06050_),
    .A1(_06051_),
    .A2(_06053_),
    .A3(_06052_),
    .S0(net497),
    .S1(net492),
    .X(_06054_));
 sky130_fd_sc_hd__o21bai_1 _12322_ (.A1(net791),
    .A2(_06054_),
    .B1_N(_06027_),
    .Y(_06055_));
 sky130_fd_sc_hd__and2_1 _12323_ (.A(_02007_),
    .B(_02076_),
    .X(_06056_));
 sky130_fd_sc_hd__inv_2 _12324_ (.A(net378),
    .Y(_06057_));
 sky130_fd_sc_hd__nor2_1 _12325_ (.A(_06041_),
    .B(net378),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _12326_ (.A(_06034_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__inv_2 _12327_ (.A(net360),
    .Y(_06060_));
 sky130_fd_sc_hd__a211o_1 _12328_ (.A1(net791),
    .A2(_06049_),
    .B1(_06055_),
    .C1(net360),
    .X(_06061_));
 sky130_fd_sc_hd__and2_1 _12329_ (.A(net719),
    .B(net380),
    .X(_06062_));
 sky130_fd_sc_hd__and2_4 _12330_ (.A(_06041_),
    .B(_06057_),
    .X(_06063_));
 sky130_fd_sc_hd__a21oi_1 _12331_ (.A1(_05989_),
    .A2(net358),
    .B1(_06062_),
    .Y(_06064_));
 sky130_fd_sc_hd__o221a_1 _12332_ (.A1(_05987_),
    .A2(_06057_),
    .B1(_06060_),
    .B2(_06064_),
    .C1(_06061_),
    .X(_06065_));
 sky130_fd_sc_hd__o2bb2a_1 _12333_ (.A1_N(_02128_),
    .A2_N(_02842_),
    .B1(_06065_),
    .B2(net478),
    .X(_06066_));
 sky130_fd_sc_hd__nor2_1 _12334_ (.A(net882),
    .B(_06066_),
    .Y(_01153_));
 sky130_fd_sc_hd__mux4_1 _12335_ (.A0(\dpath.RF.R[16][1] ),
    .A1(\dpath.RF.R[17][1] ),
    .A2(\dpath.RF.R[18][1] ),
    .A3(\dpath.RF.R[19][1] ),
    .S0(net825),
    .S1(net805),
    .X(_06067_));
 sky130_fd_sc_hd__mux4_1 _12336_ (.A0(\dpath.RF.R[20][1] ),
    .A1(net1392),
    .A2(\dpath.RF.R[22][1] ),
    .A3(\dpath.RF.R[23][1] ),
    .S0(net826),
    .S1(net806),
    .X(_06068_));
 sky130_fd_sc_hd__mux4_1 _12337_ (.A0(\dpath.RF.R[28][1] ),
    .A1(\dpath.RF.R[29][1] ),
    .A2(\dpath.RF.R[30][1] ),
    .A3(net3698),
    .S0(net825),
    .S1(net805),
    .X(_06069_));
 sky130_fd_sc_hd__mux4_1 _12338_ (.A0(\dpath.RF.R[24][1] ),
    .A1(\dpath.RF.R[25][1] ),
    .A2(\dpath.RF.R[26][1] ),
    .A3(\dpath.RF.R[27][1] ),
    .S0(net825),
    .S1(net805),
    .X(_06070_));
 sky130_fd_sc_hd__mux4_1 _12339_ (.A0(_06067_),
    .A1(_06068_),
    .A2(_06070_),
    .A3(_06069_),
    .S0(net797),
    .S1(net794),
    .X(_06071_));
 sky130_fd_sc_hd__mux4_1 _12340_ (.A0(\dpath.RF.R[0][1] ),
    .A1(\dpath.RF.R[1][1] ),
    .A2(\dpath.RF.R[2][1] ),
    .A3(\dpath.RF.R[3][1] ),
    .S0(net825),
    .S1(net805),
    .X(_06072_));
 sky130_fd_sc_hd__or2_1 _12341_ (.A(net797),
    .B(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(\dpath.RF.R[6][1] ),
    .A1(\dpath.RF.R[7][1] ),
    .S(net825),
    .X(_06074_));
 sky130_fd_sc_hd__and2_1 _12343_ (.A(net805),
    .B(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(net2548),
    .A1(net2542),
    .S(net825),
    .X(_06076_));
 sky130_fd_sc_hd__a211o_1 _12345_ (.A1(net503),
    .A2(_06076_),
    .B1(_06075_),
    .C1(net497),
    .X(_06077_));
 sky130_fd_sc_hd__mux4_1 _12346_ (.A0(\dpath.RF.R[12][1] ),
    .A1(\dpath.RF.R[13][1] ),
    .A2(\dpath.RF.R[14][1] ),
    .A3(\dpath.RF.R[15][1] ),
    .S0(net825),
    .S1(net805),
    .X(_06078_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(\dpath.RF.R[8][1] ),
    .A1(\dpath.RF.R[9][1] ),
    .S(net825),
    .X(_06079_));
 sky130_fd_sc_hd__mux2_1 _12348_ (.A0(\dpath.RF.R[10][1] ),
    .A1(\dpath.RF.R[11][1] ),
    .S(net825),
    .X(_06080_));
 sky130_fd_sc_hd__a21o_1 _12349_ (.A1(net805),
    .A2(_06080_),
    .B1(net797),
    .X(_06081_));
 sky130_fd_sc_hd__a21o_1 _12350_ (.A1(net503),
    .A2(_06079_),
    .B1(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__o211a_1 _12351_ (.A1(net497),
    .A2(_06078_),
    .B1(_06082_),
    .C1(net794),
    .X(_06083_));
 sky130_fd_sc_hd__a31o_1 _12352_ (.A1(net492),
    .A2(_06073_),
    .A3(_06077_),
    .B1(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(_06084_),
    .A1(net3699),
    .S(net791),
    .X(_06085_));
 sky130_fd_sc_hd__and2b_1 _12354_ (.A_N(_06034_),
    .B(_06058_),
    .X(_06086_));
 sky130_fd_sc_hd__and3_1 _12355_ (.A(_02007_),
    .B(_02076_),
    .C(_06022_),
    .X(_06087_));
 sky130_fd_sc_hd__a221o_1 _12356_ (.A1(_06017_),
    .A2(net358),
    .B1(_06086_),
    .B2(net716),
    .C1(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__a21oi_4 _12357_ (.A1(net364),
    .A2(_06085_),
    .B1(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__o2bb2a_1 _12358_ (.A1_N(_02123_),
    .A2_N(_02842_),
    .B1(_06089_),
    .B2(net478),
    .X(_06090_));
 sky130_fd_sc_hd__nor2_1 _12359_ (.A(net891),
    .B(_06090_),
    .Y(_01154_));
 sky130_fd_sc_hd__mux4_1 _12360_ (.A0(\dpath.RF.R[16][2] ),
    .A1(\dpath.RF.R[17][2] ),
    .A2(\dpath.RF.R[18][2] ),
    .A3(\dpath.RF.R[19][2] ),
    .S0(net827),
    .S1(net807),
    .X(_06091_));
 sky130_fd_sc_hd__mux4_1 _12361_ (.A0(\dpath.RF.R[20][2] ),
    .A1(\dpath.RF.R[21][2] ),
    .A2(\dpath.RF.R[22][2] ),
    .A3(\dpath.RF.R[23][2] ),
    .S0(net829),
    .S1(net805),
    .X(_06092_));
 sky130_fd_sc_hd__mux4_1 _12362_ (.A0(\dpath.RF.R[28][2] ),
    .A1(\dpath.RF.R[29][2] ),
    .A2(\dpath.RF.R[30][2] ),
    .A3(\dpath.RF.R[31][2] ),
    .S0(net827),
    .S1(net807),
    .X(_06093_));
 sky130_fd_sc_hd__mux4_1 _12363_ (.A0(\dpath.RF.R[24][2] ),
    .A1(\dpath.RF.R[25][2] ),
    .A2(\dpath.RF.R[26][2] ),
    .A3(\dpath.RF.R[27][2] ),
    .S0(net829),
    .S1(net805),
    .X(_06094_));
 sky130_fd_sc_hd__mux4_1 _12364_ (.A0(_06091_),
    .A1(_06092_),
    .A2(_06094_),
    .A3(_06093_),
    .S0(net797),
    .S1(net794),
    .X(_06095_));
 sky130_fd_sc_hd__mux4_1 _12365_ (.A0(\dpath.RF.R[0][2] ),
    .A1(\dpath.RF.R[1][2] ),
    .A2(\dpath.RF.R[2][2] ),
    .A3(\dpath.RF.R[3][2] ),
    .S0(net829),
    .S1(net808),
    .X(_06096_));
 sky130_fd_sc_hd__or2_1 _12366_ (.A(net797),
    .B(_06096_),
    .X(_06097_));
 sky130_fd_sc_hd__mux2_1 _12367_ (.A0(\dpath.RF.R[6][2] ),
    .A1(\dpath.RF.R[7][2] ),
    .S(net827),
    .X(_06098_));
 sky130_fd_sc_hd__and2_1 _12368_ (.A(net807),
    .B(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__mux2_1 _12369_ (.A0(\dpath.RF.R[4][2] ),
    .A1(\dpath.RF.R[5][2] ),
    .S(net827),
    .X(_06100_));
 sky130_fd_sc_hd__a211o_1 _12370_ (.A1(net503),
    .A2(_06100_),
    .B1(_06099_),
    .C1(net497),
    .X(_06101_));
 sky130_fd_sc_hd__mux4_1 _12371_ (.A0(\dpath.RF.R[12][2] ),
    .A1(\dpath.RF.R[13][2] ),
    .A2(\dpath.RF.R[14][2] ),
    .A3(\dpath.RF.R[15][2] ),
    .S0(net825),
    .S1(net805),
    .X(_06102_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(\dpath.RF.R[8][2] ),
    .A1(\dpath.RF.R[9][2] ),
    .S(net826),
    .X(_06103_));
 sky130_fd_sc_hd__mux2_1 _12373_ (.A0(\dpath.RF.R[10][2] ),
    .A1(\dpath.RF.R[11][2] ),
    .S(net826),
    .X(_06104_));
 sky130_fd_sc_hd__a21o_1 _12374_ (.A1(net806),
    .A2(_06104_),
    .B1(net797),
    .X(_06105_));
 sky130_fd_sc_hd__a21o_1 _12375_ (.A1(net503),
    .A2(_06103_),
    .B1(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__o211a_1 _12376_ (.A1(net497),
    .A2(_06102_),
    .B1(_06106_),
    .C1(net795),
    .X(_06107_));
 sky130_fd_sc_hd__a31o_1 _12377_ (.A1(net492),
    .A2(_06097_),
    .A3(_06101_),
    .B1(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(_06108_),
    .A1(_06095_),
    .S(net791),
    .X(_06109_));
 sky130_fd_sc_hd__and3_1 _12379_ (.A(_02007_),
    .B(_02076_),
    .C(_02114_),
    .X(_06110_));
 sky130_fd_sc_hd__a221o_1 _12380_ (.A1(_02099_),
    .A2(net358),
    .B1(_06086_),
    .B2(net714),
    .C1(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__a21o_1 _12381_ (.A1(net364),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__o221a_1 _12382_ (.A1(_02133_),
    .A2(_02843_),
    .B1(_06112_),
    .B2(net478),
    .C1(net862),
    .X(_01155_));
 sky130_fd_sc_hd__mux4_1 _12383_ (.A0(\dpath.RF.R[24][3] ),
    .A1(\dpath.RF.R[25][3] ),
    .A2(\dpath.RF.R[26][3] ),
    .A3(\dpath.RF.R[27][3] ),
    .S0(net819),
    .S1(net800),
    .X(_06113_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\dpath.RF.R[30][3] ),
    .A1(\dpath.RF.R[31][3] ),
    .S(net821),
    .X(_06114_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(\dpath.RF.R[28][3] ),
    .A1(\dpath.RF.R[29][3] ),
    .S(net821),
    .X(_06115_));
 sky130_fd_sc_hd__a21o_1 _12386_ (.A1(net502),
    .A2(_06115_),
    .B1(net495),
    .X(_06116_));
 sky130_fd_sc_hd__a21o_1 _12387_ (.A1(net800),
    .A2(_06114_),
    .B1(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__o211a_1 _12388_ (.A1(net796),
    .A2(_06113_),
    .B1(_06117_),
    .C1(net794),
    .X(_06118_));
 sky130_fd_sc_hd__mux4_1 _12389_ (.A0(\dpath.RF.R[20][3] ),
    .A1(\dpath.RF.R[21][3] ),
    .A2(\dpath.RF.R[22][3] ),
    .A3(\dpath.RF.R[23][3] ),
    .S0(net819),
    .S1(net800),
    .X(_06119_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(net1276),
    .A1(\dpath.RF.R[19][3] ),
    .S(net821),
    .X(_06120_));
 sky130_fd_sc_hd__mux2_1 _12391_ (.A0(\dpath.RF.R[16][3] ),
    .A1(\dpath.RF.R[17][3] ),
    .S(net821),
    .X(_06121_));
 sky130_fd_sc_hd__a21o_1 _12392_ (.A1(net502),
    .A2(_06121_),
    .B1(net796),
    .X(_06122_));
 sky130_fd_sc_hd__a21o_1 _12393_ (.A1(net800),
    .A2(_06120_),
    .B1(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__o211a_1 _12394_ (.A1(net495),
    .A2(_06119_),
    .B1(_06123_),
    .C1(net491),
    .X(_06124_));
 sky130_fd_sc_hd__or3b_1 _12395_ (.A(_06118_),
    .B(_06124_),
    .C_N(net790),
    .X(_06125_));
 sky130_fd_sc_hd__mux4_1 _12396_ (.A0(\dpath.RF.R[12][3] ),
    .A1(\dpath.RF.R[13][3] ),
    .A2(\dpath.RF.R[14][3] ),
    .A3(\dpath.RF.R[15][3] ),
    .S0(net819),
    .S1(net800),
    .X(_06126_));
 sky130_fd_sc_hd__mux4_1 _12397_ (.A0(\dpath.RF.R[8][3] ),
    .A1(\dpath.RF.R[9][3] ),
    .A2(\dpath.RF.R[10][3] ),
    .A3(\dpath.RF.R[11][3] ),
    .S0(net819),
    .S1(net800),
    .X(_06127_));
 sky130_fd_sc_hd__mux4_1 _12398_ (.A0(\dpath.RF.R[0][3] ),
    .A1(\dpath.RF.R[1][3] ),
    .A2(\dpath.RF.R[2][3] ),
    .A3(\dpath.RF.R[3][3] ),
    .S0(net819),
    .S1(net800),
    .X(_06128_));
 sky130_fd_sc_hd__mux4_1 _12399_ (.A0(\dpath.RF.R[4][3] ),
    .A1(\dpath.RF.R[5][3] ),
    .A2(\dpath.RF.R[6][3] ),
    .A3(\dpath.RF.R[7][3] ),
    .S0(net819),
    .S1(net800),
    .X(_06129_));
 sky130_fd_sc_hd__mux4_1 _12400_ (.A0(_06126_),
    .A1(_06127_),
    .A2(_06129_),
    .A3(_06128_),
    .S0(net495),
    .S1(net491),
    .X(_06130_));
 sky130_fd_sc_hd__or2_1 _12401_ (.A(net790),
    .B(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__and3_1 _12402_ (.A(net364),
    .B(_06125_),
    .C(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__a22o_1 _12403_ (.A1(net713),
    .A2(net380),
    .B1(net358),
    .B2(_02163_),
    .X(_06133_));
 sky130_fd_sc_hd__a21o_1 _12404_ (.A1(_02183_),
    .A2(net378),
    .B1(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__a21oi_4 _12405_ (.A1(net360),
    .A2(_06134_),
    .B1(_06132_),
    .Y(_06135_));
 sky130_fd_sc_hd__o2bb2a_1 _12406_ (.A1_N(_02187_),
    .A2_N(_02842_),
    .B1(_06135_),
    .B2(net478),
    .X(_06136_));
 sky130_fd_sc_hd__nor2_1 _12407_ (.A(net890),
    .B(_06136_),
    .Y(_01156_));
 sky130_fd_sc_hd__mux4_1 _12408_ (.A0(net2538),
    .A1(\dpath.RF.R[25][4] ),
    .A2(net1566),
    .A3(net2776),
    .S0(net820),
    .S1(net801),
    .X(_06137_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(net1706),
    .A1(net2458),
    .S(net820),
    .X(_06138_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(\dpath.RF.R[28][4] ),
    .A1(\dpath.RF.R[29][4] ),
    .S(net820),
    .X(_06139_));
 sky130_fd_sc_hd__a21o_1 _12411_ (.A1(net502),
    .A2(_06139_),
    .B1(net495),
    .X(_06140_));
 sky130_fd_sc_hd__a21o_1 _12412_ (.A1(net804),
    .A2(_06138_),
    .B1(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__o211a_1 _12413_ (.A1(net796),
    .A2(_06137_),
    .B1(_06141_),
    .C1(net794),
    .X(_06142_));
 sky130_fd_sc_hd__mux4_1 _12414_ (.A0(\dpath.RF.R[20][4] ),
    .A1(\dpath.RF.R[21][4] ),
    .A2(\dpath.RF.R[22][4] ),
    .A3(net2526),
    .S0(net820),
    .S1(net801),
    .X(_06143_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(\dpath.RF.R[18][4] ),
    .A1(\dpath.RF.R[19][4] ),
    .S(net821),
    .X(_06144_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(\dpath.RF.R[16][4] ),
    .A1(\dpath.RF.R[17][4] ),
    .S(net820),
    .X(_06145_));
 sky130_fd_sc_hd__a21o_1 _12417_ (.A1(net502),
    .A2(_06145_),
    .B1(net796),
    .X(_06146_));
 sky130_fd_sc_hd__a21o_1 _12418_ (.A1(net801),
    .A2(_06144_),
    .B1(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__o211a_1 _12419_ (.A1(net495),
    .A2(_06143_),
    .B1(_06147_),
    .C1(net491),
    .X(_06148_));
 sky130_fd_sc_hd__or3b_1 _12420_ (.A(_06142_),
    .B(_06148_),
    .C_N(net790),
    .X(_06149_));
 sky130_fd_sc_hd__mux4_1 _12421_ (.A0(\dpath.RF.R[12][4] ),
    .A1(\dpath.RF.R[13][4] ),
    .A2(\dpath.RF.R[14][4] ),
    .A3(\dpath.RF.R[15][4] ),
    .S0(net820),
    .S1(net801),
    .X(_06150_));
 sky130_fd_sc_hd__mux4_1 _12422_ (.A0(\dpath.RF.R[8][4] ),
    .A1(\dpath.RF.R[9][4] ),
    .A2(\dpath.RF.R[10][4] ),
    .A3(\dpath.RF.R[11][4] ),
    .S0(net820),
    .S1(net801),
    .X(_06151_));
 sky130_fd_sc_hd__mux4_1 _12423_ (.A0(\dpath.RF.R[0][4] ),
    .A1(\dpath.RF.R[1][4] ),
    .A2(\dpath.RF.R[2][4] ),
    .A3(\dpath.RF.R[3][4] ),
    .S0(net820),
    .S1(net801),
    .X(_06152_));
 sky130_fd_sc_hd__mux4_1 _12424_ (.A0(\dpath.RF.R[4][4] ),
    .A1(\dpath.RF.R[5][4] ),
    .A2(\dpath.RF.R[6][4] ),
    .A3(\dpath.RF.R[7][4] ),
    .S0(net820),
    .S1(net801),
    .X(_06153_));
 sky130_fd_sc_hd__mux4_1 _12425_ (.A0(_06150_),
    .A1(_06151_),
    .A2(_06153_),
    .A3(_06152_),
    .S0(net495),
    .S1(net491),
    .X(_06154_));
 sky130_fd_sc_hd__or2_1 _12426_ (.A(net790),
    .B(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__and3_1 _12427_ (.A(net364),
    .B(_06149_),
    .C(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__a22o_1 _12428_ (.A1(net3267),
    .A2(net380),
    .B1(net358),
    .B2(_02217_),
    .X(_06157_));
 sky130_fd_sc_hd__a21o_1 _12429_ (.A1(_02246_),
    .A2(net378),
    .B1(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__a21oi_4 _12430_ (.A1(net360),
    .A2(_06158_),
    .B1(_06156_),
    .Y(_06159_));
 sky130_fd_sc_hd__o2bb2a_1 _12431_ (.A1_N(_02250_),
    .A2_N(_02842_),
    .B1(_06159_),
    .B2(net478),
    .X(_06160_));
 sky130_fd_sc_hd__nor2_1 _12432_ (.A(net890),
    .B(_06160_),
    .Y(_01157_));
 sky130_fd_sc_hd__mux4_1 _12433_ (.A0(net2424),
    .A1(net3134),
    .A2(net2110),
    .A3(net2062),
    .S0(net823),
    .S1(net803),
    .X(_06161_));
 sky130_fd_sc_hd__mux2_1 _12434_ (.A0(net1556),
    .A1(net3104),
    .S(net823),
    .X(_06162_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(\dpath.RF.R[28][5] ),
    .A1(\dpath.RF.R[29][5] ),
    .S(net823),
    .X(_06163_));
 sky130_fd_sc_hd__a21o_1 _12436_ (.A1(net502),
    .A2(_06163_),
    .B1(net496),
    .X(_06164_));
 sky130_fd_sc_hd__a21o_1 _12437_ (.A1(net803),
    .A2(_06162_),
    .B1(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__o211a_1 _12438_ (.A1(net796),
    .A2(_06161_),
    .B1(_06165_),
    .C1(net794),
    .X(_06166_));
 sky130_fd_sc_hd__mux4_1 _12439_ (.A0(net1398),
    .A1(net2590),
    .A2(net2574),
    .A3(net2036),
    .S0(net821),
    .S1(net801),
    .X(_06167_));
 sky130_fd_sc_hd__mux2_1 _12440_ (.A0(net2186),
    .A1(net2008),
    .S(net823),
    .X(_06168_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(\dpath.RF.R[16][5] ),
    .A1(\dpath.RF.R[17][5] ),
    .S(net823),
    .X(_06169_));
 sky130_fd_sc_hd__a21o_1 _12442_ (.A1(net502),
    .A2(_06169_),
    .B1(net796),
    .X(_06170_));
 sky130_fd_sc_hd__a21o_1 _12443_ (.A1(net801),
    .A2(_06168_),
    .B1(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__o211a_1 _12444_ (.A1(net495),
    .A2(_06167_),
    .B1(_06171_),
    .C1(net491),
    .X(_06172_));
 sky130_fd_sc_hd__or3b_1 _12445_ (.A(_06166_),
    .B(_06172_),
    .C_N(net790),
    .X(_06173_));
 sky130_fd_sc_hd__mux4_1 _12446_ (.A0(\dpath.RF.R[12][5] ),
    .A1(\dpath.RF.R[13][5] ),
    .A2(\dpath.RF.R[14][5] ),
    .A3(\dpath.RF.R[15][5] ),
    .S0(net823),
    .S1(net803),
    .X(_06174_));
 sky130_fd_sc_hd__mux4_1 _12447_ (.A0(\dpath.RF.R[8][5] ),
    .A1(\dpath.RF.R[9][5] ),
    .A2(\dpath.RF.R[10][5] ),
    .A3(\dpath.RF.R[11][5] ),
    .S0(net823),
    .S1(net803),
    .X(_06175_));
 sky130_fd_sc_hd__mux4_1 _12448_ (.A0(\dpath.RF.R[0][5] ),
    .A1(\dpath.RF.R[1][5] ),
    .A2(\dpath.RF.R[2][5] ),
    .A3(\dpath.RF.R[3][5] ),
    .S0(net821),
    .S1(net801),
    .X(_06176_));
 sky130_fd_sc_hd__mux4_1 _12449_ (.A0(\dpath.RF.R[4][5] ),
    .A1(\dpath.RF.R[5][5] ),
    .A2(\dpath.RF.R[6][5] ),
    .A3(\dpath.RF.R[7][5] ),
    .S0(net821),
    .S1(net804),
    .X(_06177_));
 sky130_fd_sc_hd__mux4_1 _12450_ (.A0(_06174_),
    .A1(_06175_),
    .A2(_06177_),
    .A3(_06176_),
    .S0(net495),
    .S1(net491),
    .X(_06178_));
 sky130_fd_sc_hd__or2_1 _12451_ (.A(net790),
    .B(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__and3_1 _12452_ (.A(net364),
    .B(_06173_),
    .C(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__a22o_1 _12453_ (.A1(net708),
    .A2(net380),
    .B1(net358),
    .B2(_02284_),
    .X(_06181_));
 sky130_fd_sc_hd__a21o_1 _12454_ (.A1(_02316_),
    .A2(net378),
    .B1(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__a21oi_4 _12455_ (.A1(net360),
    .A2(net3625),
    .B1(_06180_),
    .Y(_06183_));
 sky130_fd_sc_hd__o2bb2a_1 _12456_ (.A1_N(net3392),
    .A2_N(_02842_),
    .B1(_06183_),
    .B2(net478),
    .X(_06184_));
 sky130_fd_sc_hd__nor2_1 _12457_ (.A(net891),
    .B(_06184_),
    .Y(_01158_));
 sky130_fd_sc_hd__mux4_1 _12458_ (.A0(net1536),
    .A1(net2902),
    .A2(\dpath.RF.R[26][6] ),
    .A3(net2340),
    .S0(net820),
    .S1(net801),
    .X(_06185_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(net1942),
    .A1(net3042),
    .S(net820),
    .X(_06186_));
 sky130_fd_sc_hd__mux2_1 _12460_ (.A0(\dpath.RF.R[28][6] ),
    .A1(\dpath.RF.R[29][6] ),
    .S(net821),
    .X(_06187_));
 sky130_fd_sc_hd__a21o_1 _12461_ (.A1(net502),
    .A2(_06187_),
    .B1(net495),
    .X(_06188_));
 sky130_fd_sc_hd__a21o_1 _12462_ (.A1(net804),
    .A2(_06186_),
    .B1(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__o211a_1 _12463_ (.A1(net796),
    .A2(_06185_),
    .B1(_06189_),
    .C1(net794),
    .X(_06190_));
 sky130_fd_sc_hd__mux4_1 _12464_ (.A0(net2454),
    .A1(net3697),
    .A2(\dpath.RF.R[22][6] ),
    .A3(net3136),
    .S0(net820),
    .S1(net801),
    .X(_06191_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(net2630),
    .A1(net2426),
    .S(net825),
    .X(_06192_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(\dpath.RF.R[16][6] ),
    .A1(\dpath.RF.R[17][6] ),
    .S(net825),
    .X(_06193_));
 sky130_fd_sc_hd__a21o_1 _12467_ (.A1(net502),
    .A2(_06193_),
    .B1(net796),
    .X(_06194_));
 sky130_fd_sc_hd__a21o_1 _12468_ (.A1(net805),
    .A2(_06192_),
    .B1(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__o211a_1 _12469_ (.A1(net495),
    .A2(_06191_),
    .B1(_06195_),
    .C1(net491),
    .X(_06196_));
 sky130_fd_sc_hd__or3b_1 _12470_ (.A(_06190_),
    .B(_06196_),
    .C_N(net790),
    .X(_06197_));
 sky130_fd_sc_hd__mux4_1 _12471_ (.A0(\dpath.RF.R[12][6] ),
    .A1(\dpath.RF.R[13][6] ),
    .A2(\dpath.RF.R[14][6] ),
    .A3(\dpath.RF.R[15][6] ),
    .S0(net820),
    .S1(net801),
    .X(_06198_));
 sky130_fd_sc_hd__mux4_1 _12472_ (.A0(\dpath.RF.R[8][6] ),
    .A1(\dpath.RF.R[9][6] ),
    .A2(\dpath.RF.R[10][6] ),
    .A3(\dpath.RF.R[11][6] ),
    .S0(net820),
    .S1(net801),
    .X(_06199_));
 sky130_fd_sc_hd__mux4_1 _12473_ (.A0(\dpath.RF.R[0][6] ),
    .A1(\dpath.RF.R[1][6] ),
    .A2(\dpath.RF.R[2][6] ),
    .A3(\dpath.RF.R[3][6] ),
    .S0(net820),
    .S1(net801),
    .X(_06200_));
 sky130_fd_sc_hd__mux4_1 _12474_ (.A0(\dpath.RF.R[4][6] ),
    .A1(\dpath.RF.R[5][6] ),
    .A2(\dpath.RF.R[6][6] ),
    .A3(\dpath.RF.R[7][6] ),
    .S0(net820),
    .S1(net801),
    .X(_06201_));
 sky130_fd_sc_hd__mux4_1 _12475_ (.A0(_06198_),
    .A1(_06199_),
    .A2(_06201_),
    .A3(_06200_),
    .S0(net495),
    .S1(net491),
    .X(_06202_));
 sky130_fd_sc_hd__or2_1 _12476_ (.A(net790),
    .B(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__and3_1 _12477_ (.A(net364),
    .B(_06197_),
    .C(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__a22o_1 _12478_ (.A1(net707),
    .A2(net380),
    .B1(net358),
    .B2(_02347_),
    .X(_06205_));
 sky130_fd_sc_hd__a21o_1 _12479_ (.A1(_02387_),
    .A2(net378),
    .B1(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__a21oi_4 _12480_ (.A1(net360),
    .A2(_06206_),
    .B1(_06204_),
    .Y(_06207_));
 sky130_fd_sc_hd__o2bb2a_1 _12481_ (.A1_N(net3452),
    .A2_N(_02125_),
    .B1(_06207_),
    .B2(net478),
    .X(_06208_));
 sky130_fd_sc_hd__nor2_1 _12482_ (.A(net890),
    .B(_06208_),
    .Y(_01159_));
 sky130_fd_sc_hd__mux4_1 _12483_ (.A0(\dpath.RF.R[24][7] ),
    .A1(\dpath.RF.R[25][7] ),
    .A2(\dpath.RF.R[26][7] ),
    .A3(\dpath.RF.R[27][7] ),
    .S0(net819),
    .S1(net800),
    .X(_06209_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(\dpath.RF.R[30][7] ),
    .A1(\dpath.RF.R[31][7] ),
    .S(net819),
    .X(_06210_));
 sky130_fd_sc_hd__mux2_1 _12485_ (.A0(\dpath.RF.R[28][7] ),
    .A1(\dpath.RF.R[29][7] ),
    .S(net819),
    .X(_06211_));
 sky130_fd_sc_hd__a21o_1 _12486_ (.A1(net502),
    .A2(_06211_),
    .B1(net495),
    .X(_06212_));
 sky130_fd_sc_hd__a21o_1 _12487_ (.A1(net800),
    .A2(_06210_),
    .B1(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__o211a_1 _12488_ (.A1(net796),
    .A2(_06209_),
    .B1(_06213_),
    .C1(net794),
    .X(_06214_));
 sky130_fd_sc_hd__mux4_1 _12489_ (.A0(\dpath.RF.R[20][7] ),
    .A1(\dpath.RF.R[21][7] ),
    .A2(\dpath.RF.R[22][7] ),
    .A3(\dpath.RF.R[23][7] ),
    .S0(net819),
    .S1(net800),
    .X(_06215_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(net1336),
    .A1(\dpath.RF.R[19][7] ),
    .S(net819),
    .X(_06216_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(\dpath.RF.R[16][7] ),
    .A1(\dpath.RF.R[17][7] ),
    .S(net819),
    .X(_06217_));
 sky130_fd_sc_hd__a21o_1 _12492_ (.A1(net502),
    .A2(_06217_),
    .B1(net796),
    .X(_06218_));
 sky130_fd_sc_hd__a21o_1 _12493_ (.A1(net800),
    .A2(_06216_),
    .B1(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__o211a_1 _12494_ (.A1(net495),
    .A2(_06215_),
    .B1(_06219_),
    .C1(net491),
    .X(_06220_));
 sky130_fd_sc_hd__or3b_1 _12495_ (.A(_06214_),
    .B(_06220_),
    .C_N(net790),
    .X(_06221_));
 sky130_fd_sc_hd__mux4_1 _12496_ (.A0(\dpath.RF.R[12][7] ),
    .A1(\dpath.RF.R[13][7] ),
    .A2(\dpath.RF.R[14][7] ),
    .A3(\dpath.RF.R[15][7] ),
    .S0(net819),
    .S1(net800),
    .X(_06222_));
 sky130_fd_sc_hd__mux4_1 _12497_ (.A0(\dpath.RF.R[8][7] ),
    .A1(\dpath.RF.R[9][7] ),
    .A2(\dpath.RF.R[10][7] ),
    .A3(\dpath.RF.R[11][7] ),
    .S0(net821),
    .S1(net804),
    .X(_06223_));
 sky130_fd_sc_hd__mux4_1 _12498_ (.A0(\dpath.RF.R[0][7] ),
    .A1(\dpath.RF.R[1][7] ),
    .A2(\dpath.RF.R[2][7] ),
    .A3(\dpath.RF.R[3][7] ),
    .S0(net819),
    .S1(net800),
    .X(_06224_));
 sky130_fd_sc_hd__mux4_1 _12499_ (.A0(\dpath.RF.R[4][7] ),
    .A1(\dpath.RF.R[5][7] ),
    .A2(\dpath.RF.R[6][7] ),
    .A3(\dpath.RF.R[7][7] ),
    .S0(net821),
    .S1(net804),
    .X(_06225_));
 sky130_fd_sc_hd__mux4_1 _12500_ (.A0(_06222_),
    .A1(_06223_),
    .A2(_06225_),
    .A3(_06224_),
    .S0(net495),
    .S1(net491),
    .X(_06226_));
 sky130_fd_sc_hd__or2_1 _12501_ (.A(net790),
    .B(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__and3_1 _12502_ (.A(net364),
    .B(_06221_),
    .C(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__a22o_1 _12503_ (.A1(net704),
    .A2(net380),
    .B1(net358),
    .B2(_02418_),
    .X(_06229_));
 sky130_fd_sc_hd__a21o_1 _12504_ (.A1(_02459_),
    .A2(net378),
    .B1(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__a21oi_4 _12505_ (.A1(net360),
    .A2(_06230_),
    .B1(_06228_),
    .Y(_06231_));
 sky130_fd_sc_hd__o2bb2a_1 _12506_ (.A1_N(net3420),
    .A2_N(_02842_),
    .B1(_06231_),
    .B2(net478),
    .X(_06232_));
 sky130_fd_sc_hd__nor2_1 _12507_ (.A(net891),
    .B(_06232_),
    .Y(_01160_));
 sky130_fd_sc_hd__mux4_1 _12508_ (.A0(\dpath.RF.R[24][8] ),
    .A1(\dpath.RF.R[25][8] ),
    .A2(\dpath.RF.R[26][8] ),
    .A3(\dpath.RF.R[27][8] ),
    .S0(net827),
    .S1(net807),
    .X(_06233_));
 sky130_fd_sc_hd__mux2_1 _12509_ (.A0(\dpath.RF.R[30][8] ),
    .A1(\dpath.RF.R[31][8] ),
    .S(net827),
    .X(_06234_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(\dpath.RF.R[28][8] ),
    .A1(\dpath.RF.R[29][8] ),
    .S(net828),
    .X(_06235_));
 sky130_fd_sc_hd__a21o_1 _12511_ (.A1(net503),
    .A2(_06235_),
    .B1(net497),
    .X(_06236_));
 sky130_fd_sc_hd__a21o_1 _12512_ (.A1(net807),
    .A2(_06234_),
    .B1(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__o211a_1 _12513_ (.A1(net797),
    .A2(_06233_),
    .B1(_06237_),
    .C1(net795),
    .X(_06238_));
 sky130_fd_sc_hd__mux4_1 _12514_ (.A0(\dpath.RF.R[20][8] ),
    .A1(\dpath.RF.R[21][8] ),
    .A2(\dpath.RF.R[22][8] ),
    .A3(\dpath.RF.R[23][8] ),
    .S0(net827),
    .S1(net807),
    .X(_06239_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(\dpath.RF.R[18][8] ),
    .A1(\dpath.RF.R[19][8] ),
    .S(net828),
    .X(_06240_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(\dpath.RF.R[16][8] ),
    .A1(\dpath.RF.R[17][8] ),
    .S(net828),
    .X(_06241_));
 sky130_fd_sc_hd__a21o_1 _12517_ (.A1(net503),
    .A2(_06241_),
    .B1(_00002_),
    .X(_06242_));
 sky130_fd_sc_hd__a21o_1 _12518_ (.A1(net807),
    .A2(_06240_),
    .B1(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__o211a_1 _12519_ (.A1(net497),
    .A2(_06239_),
    .B1(_06243_),
    .C1(net492),
    .X(_06244_));
 sky130_fd_sc_hd__or3b_1 _12520_ (.A(_06238_),
    .B(_06244_),
    .C_N(net791),
    .X(_06245_));
 sky130_fd_sc_hd__mux4_1 _12521_ (.A0(\dpath.RF.R[12][8] ),
    .A1(\dpath.RF.R[13][8] ),
    .A2(\dpath.RF.R[14][8] ),
    .A3(\dpath.RF.R[15][8] ),
    .S0(net828),
    .S1(net807),
    .X(_06246_));
 sky130_fd_sc_hd__mux4_1 _12522_ (.A0(\dpath.RF.R[8][8] ),
    .A1(\dpath.RF.R[9][8] ),
    .A2(\dpath.RF.R[10][8] ),
    .A3(\dpath.RF.R[11][8] ),
    .S0(net826),
    .S1(net806),
    .X(_06247_));
 sky130_fd_sc_hd__mux4_1 _12523_ (.A0(\dpath.RF.R[0][8] ),
    .A1(\dpath.RF.R[1][8] ),
    .A2(\dpath.RF.R[2][8] ),
    .A3(\dpath.RF.R[3][8] ),
    .S0(net827),
    .S1(net807),
    .X(_06248_));
 sky130_fd_sc_hd__mux4_1 _12524_ (.A0(\dpath.RF.R[4][8] ),
    .A1(\dpath.RF.R[5][8] ),
    .A2(\dpath.RF.R[6][8] ),
    .A3(\dpath.RF.R[7][8] ),
    .S0(net827),
    .S1(net807),
    .X(_06249_));
 sky130_fd_sc_hd__mux4_1 _12525_ (.A0(_06246_),
    .A1(_06247_),
    .A2(_06249_),
    .A3(_06248_),
    .S0(net497),
    .S1(net492),
    .X(_06250_));
 sky130_fd_sc_hd__or2_1 _12526_ (.A(net791),
    .B(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__and3_1 _12527_ (.A(net364),
    .B(_06245_),
    .C(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__a22o_1 _12528_ (.A1(net703),
    .A2(net380),
    .B1(net358),
    .B2(_02496_),
    .X(_06253_));
 sky130_fd_sc_hd__a21o_1 _12529_ (.A1(_02551_),
    .A2(net378),
    .B1(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__a21oi_2 _12530_ (.A1(net360),
    .A2(_06254_),
    .B1(_06252_),
    .Y(_06255_));
 sky130_fd_sc_hd__o2bb2a_1 _12531_ (.A1_N(net3421),
    .A2_N(_02842_),
    .B1(_06255_),
    .B2(net478),
    .X(_06256_));
 sky130_fd_sc_hd__nor2_1 _12532_ (.A(net891),
    .B(_06256_),
    .Y(_01161_));
 sky130_fd_sc_hd__mux4_1 _12533_ (.A0(net1606),
    .A1(net1644),
    .A2(net1474),
    .A3(net2416),
    .S0(net826),
    .S1(net806),
    .X(_06257_));
 sky130_fd_sc_hd__mux2_1 _12534_ (.A0(net2164),
    .A1(net2958),
    .S(net828),
    .X(_06258_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(\dpath.RF.R[28][9] ),
    .A1(\dpath.RF.R[29][9] ),
    .S(net828),
    .X(_06259_));
 sky130_fd_sc_hd__a21o_1 _12536_ (.A1(net503),
    .A2(_06259_),
    .B1(net497),
    .X(_06260_));
 sky130_fd_sc_hd__a21o_1 _12537_ (.A1(net806),
    .A2(_06258_),
    .B1(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__o211a_1 _12538_ (.A1(net797),
    .A2(_06257_),
    .B1(_06261_),
    .C1(net795),
    .X(_06262_));
 sky130_fd_sc_hd__mux4_1 _12539_ (.A0(net2056),
    .A1(net1472),
    .A2(net3703),
    .A3(net3004),
    .S0(net826),
    .S1(net806),
    .X(_06263_));
 sky130_fd_sc_hd__mux2_1 _12540_ (.A0(net1820),
    .A1(net2348),
    .S(net826),
    .X(_06264_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\dpath.RF.R[16][9] ),
    .A1(\dpath.RF.R[17][9] ),
    .S(net826),
    .X(_06265_));
 sky130_fd_sc_hd__a21o_1 _12542_ (.A1(net503),
    .A2(_06265_),
    .B1(_00002_),
    .X(_06266_));
 sky130_fd_sc_hd__a21o_1 _12543_ (.A1(net806),
    .A2(_06264_),
    .B1(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__o211a_1 _12544_ (.A1(_01789_),
    .A2(_06263_),
    .B1(_06267_),
    .C1(net492),
    .X(_06268_));
 sky130_fd_sc_hd__or3b_1 _12545_ (.A(_06262_),
    .B(_06268_),
    .C_N(net791),
    .X(_06269_));
 sky130_fd_sc_hd__mux4_1 _12546_ (.A0(\dpath.RF.R[12][9] ),
    .A1(\dpath.RF.R[13][9] ),
    .A2(\dpath.RF.R[14][9] ),
    .A3(\dpath.RF.R[15][9] ),
    .S0(net826),
    .S1(net806),
    .X(_06270_));
 sky130_fd_sc_hd__mux4_1 _12547_ (.A0(\dpath.RF.R[8][9] ),
    .A1(\dpath.RF.R[9][9] ),
    .A2(\dpath.RF.R[10][9] ),
    .A3(\dpath.RF.R[11][9] ),
    .S0(net823),
    .S1(net803),
    .X(_06271_));
 sky130_fd_sc_hd__mux4_1 _12548_ (.A0(\dpath.RF.R[0][9] ),
    .A1(\dpath.RF.R[1][9] ),
    .A2(\dpath.RF.R[2][9] ),
    .A3(\dpath.RF.R[3][9] ),
    .S0(net826),
    .S1(net806),
    .X(_06272_));
 sky130_fd_sc_hd__mux4_1 _12549_ (.A0(\dpath.RF.R[4][9] ),
    .A1(\dpath.RF.R[5][9] ),
    .A2(\dpath.RF.R[6][9] ),
    .A3(\dpath.RF.R[7][9] ),
    .S0(net826),
    .S1(net806),
    .X(_06273_));
 sky130_fd_sc_hd__mux4_1 _12550_ (.A0(_06270_),
    .A1(_06271_),
    .A2(_06273_),
    .A3(_06272_),
    .S0(_01789_),
    .S1(net492),
    .X(_06274_));
 sky130_fd_sc_hd__or2_1 _12551_ (.A(net791),
    .B(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__and3_1 _12552_ (.A(net364),
    .B(_06269_),
    .C(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__a22o_1 _12553_ (.A1(net700),
    .A2(net380),
    .B1(net358),
    .B2(_02584_),
    .X(_06277_));
 sky130_fd_sc_hd__a21o_1 _12554_ (.A1(_02640_),
    .A2(net378),
    .B1(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__a21oi_4 _12555_ (.A1(net360),
    .A2(_06278_),
    .B1(_06276_),
    .Y(_06279_));
 sky130_fd_sc_hd__o2bb2a_1 _12556_ (.A1_N(net3461),
    .A2_N(_02842_),
    .B1(_06279_),
    .B2(net478),
    .X(_06280_));
 sky130_fd_sc_hd__nor2_1 _12557_ (.A(net891),
    .B(_06280_),
    .Y(_01162_));
 sky130_fd_sc_hd__mux4_1 _12558_ (.A0(net1094),
    .A1(net2878),
    .A2(net1324),
    .A3(net3694),
    .S0(net827),
    .S1(net807),
    .X(_06281_));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(net1660),
    .A1(net2624),
    .S(net827),
    .X(_06282_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(\dpath.RF.R[28][10] ),
    .A1(\dpath.RF.R[29][10] ),
    .S(net828),
    .X(_06283_));
 sky130_fd_sc_hd__a21o_1 _12561_ (.A1(net503),
    .A2(_06283_),
    .B1(net497),
    .X(_06284_));
 sky130_fd_sc_hd__a21o_1 _12562_ (.A1(net807),
    .A2(_06282_),
    .B1(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__o211a_1 _12563_ (.A1(net797),
    .A2(_06281_),
    .B1(_06285_),
    .C1(net794),
    .X(_06286_));
 sky130_fd_sc_hd__mux4_1 _12564_ (.A0(net1716),
    .A1(net1944),
    .A2(net1794),
    .A3(net2118),
    .S0(net827),
    .S1(net807),
    .X(_06287_));
 sky130_fd_sc_hd__mux2_1 _12565_ (.A0(net1854),
    .A1(net1456),
    .S(net827),
    .X(_06288_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\dpath.RF.R[16][10] ),
    .A1(\dpath.RF.R[17][10] ),
    .S(net827),
    .X(_06289_));
 sky130_fd_sc_hd__a21o_1 _12567_ (.A1(net503),
    .A2(_06289_),
    .B1(net797),
    .X(_06290_));
 sky130_fd_sc_hd__a21o_1 _12568_ (.A1(net807),
    .A2(_06288_),
    .B1(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__o211a_1 _12569_ (.A1(net497),
    .A2(_06287_),
    .B1(_06291_),
    .C1(net492),
    .X(_06292_));
 sky130_fd_sc_hd__or3b_1 _12570_ (.A(_06286_),
    .B(_06292_),
    .C_N(net791),
    .X(_06293_));
 sky130_fd_sc_hd__mux4_1 _12571_ (.A0(\dpath.RF.R[12][10] ),
    .A1(\dpath.RF.R[13][10] ),
    .A2(\dpath.RF.R[14][10] ),
    .A3(\dpath.RF.R[15][10] ),
    .S0(net827),
    .S1(net807),
    .X(_06294_));
 sky130_fd_sc_hd__mux4_1 _12572_ (.A0(\dpath.RF.R[8][10] ),
    .A1(\dpath.RF.R[9][10] ),
    .A2(\dpath.RF.R[10][10] ),
    .A3(\dpath.RF.R[11][10] ),
    .S0(net826),
    .S1(net806),
    .X(_06295_));
 sky130_fd_sc_hd__mux4_1 _12573_ (.A0(\dpath.RF.R[0][10] ),
    .A1(\dpath.RF.R[1][10] ),
    .A2(\dpath.RF.R[2][10] ),
    .A3(\dpath.RF.R[3][10] ),
    .S0(net827),
    .S1(net807),
    .X(_06296_));
 sky130_fd_sc_hd__mux4_1 _12574_ (.A0(\dpath.RF.R[4][10] ),
    .A1(\dpath.RF.R[5][10] ),
    .A2(\dpath.RF.R[6][10] ),
    .A3(\dpath.RF.R[7][10] ),
    .S0(net826),
    .S1(net806),
    .X(_06297_));
 sky130_fd_sc_hd__mux4_1 _12575_ (.A0(_06294_),
    .A1(_06295_),
    .A2(_06297_),
    .A3(_06296_),
    .S0(net497),
    .S1(net492),
    .X(_06298_));
 sky130_fd_sc_hd__or2_1 _12576_ (.A(net791),
    .B(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__and3_1 _12577_ (.A(net364),
    .B(_06293_),
    .C(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__a22o_1 _12578_ (.A1(net698),
    .A2(net380),
    .B1(net358),
    .B2(_02674_),
    .X(_06301_));
 sky130_fd_sc_hd__a21o_1 _12579_ (.A1(_02740_),
    .A2(net378),
    .B1(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__a21oi_2 _12580_ (.A1(net360),
    .A2(_06302_),
    .B1(_06300_),
    .Y(_06303_));
 sky130_fd_sc_hd__o2bb2a_1 _12581_ (.A1_N(net3435),
    .A2_N(_02842_),
    .B1(_06303_),
    .B2(net478),
    .X(_06304_));
 sky130_fd_sc_hd__nor2_1 _12582_ (.A(net891),
    .B(_06304_),
    .Y(_01163_));
 sky130_fd_sc_hd__mux4_1 _12583_ (.A0(\dpath.RF.R[24][11] ),
    .A1(\dpath.RF.R[25][11] ),
    .A2(\dpath.RF.R[26][11] ),
    .A3(\dpath.RF.R[27][11] ),
    .S0(net822),
    .S1(net802),
    .X(_06305_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(\dpath.RF.R[30][11] ),
    .A1(\dpath.RF.R[31][11] ),
    .S(net822),
    .X(_06306_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(\dpath.RF.R[28][11] ),
    .A1(\dpath.RF.R[29][11] ),
    .S(net822),
    .X(_06307_));
 sky130_fd_sc_hd__a21o_1 _12586_ (.A1(net502),
    .A2(_06307_),
    .B1(net496),
    .X(_06308_));
 sky130_fd_sc_hd__a21o_1 _12587_ (.A1(net802),
    .A2(_06306_),
    .B1(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__o211a_1 _12588_ (.A1(net796),
    .A2(_06305_),
    .B1(_06309_),
    .C1(net794),
    .X(_06310_));
 sky130_fd_sc_hd__mux4_1 _12589_ (.A0(\dpath.RF.R[20][11] ),
    .A1(\dpath.RF.R[21][11] ),
    .A2(\dpath.RF.R[22][11] ),
    .A3(\dpath.RF.R[23][11] ),
    .S0(net822),
    .S1(net802),
    .X(_06311_));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(\dpath.RF.R[18][11] ),
    .A1(\dpath.RF.R[19][11] ),
    .S(net822),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(\dpath.RF.R[16][11] ),
    .A1(\dpath.RF.R[17][11] ),
    .S(net822),
    .X(_06313_));
 sky130_fd_sc_hd__a21o_1 _12592_ (.A1(net502),
    .A2(_06313_),
    .B1(net796),
    .X(_06314_));
 sky130_fd_sc_hd__a21o_1 _12593_ (.A1(net802),
    .A2(_06312_),
    .B1(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__o211a_1 _12594_ (.A1(net496),
    .A2(_06311_),
    .B1(_06315_),
    .C1(net492),
    .X(_06316_));
 sky130_fd_sc_hd__or3b_1 _12595_ (.A(_06310_),
    .B(_06316_),
    .C_N(net790),
    .X(_06317_));
 sky130_fd_sc_hd__mux4_1 _12596_ (.A0(\dpath.RF.R[12][11] ),
    .A1(\dpath.RF.R[13][11] ),
    .A2(\dpath.RF.R[14][11] ),
    .A3(\dpath.RF.R[15][11] ),
    .S0(net822),
    .S1(net802),
    .X(_06318_));
 sky130_fd_sc_hd__mux4_1 _12597_ (.A0(\dpath.RF.R[8][11] ),
    .A1(\dpath.RF.R[9][11] ),
    .A2(\dpath.RF.R[10][11] ),
    .A3(\dpath.RF.R[11][11] ),
    .S0(net822),
    .S1(net802),
    .X(_06319_));
 sky130_fd_sc_hd__mux4_1 _12598_ (.A0(\dpath.RF.R[0][11] ),
    .A1(\dpath.RF.R[1][11] ),
    .A2(\dpath.RF.R[2][11] ),
    .A3(\dpath.RF.R[3][11] ),
    .S0(net819),
    .S1(net800),
    .X(_06320_));
 sky130_fd_sc_hd__mux4_1 _12599_ (.A0(\dpath.RF.R[4][11] ),
    .A1(\dpath.RF.R[5][11] ),
    .A2(\dpath.RF.R[6][11] ),
    .A3(\dpath.RF.R[7][11] ),
    .S0(net819),
    .S1(net800),
    .X(_06321_));
 sky130_fd_sc_hd__mux4_1 _12600_ (.A0(_06318_),
    .A1(_06319_),
    .A2(_06321_),
    .A3(_06320_),
    .S0(net495),
    .S1(net491),
    .X(_06322_));
 sky130_fd_sc_hd__or2_1 _12601_ (.A(net791),
    .B(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__and3_1 _12602_ (.A(net364),
    .B(_06317_),
    .C(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__a22o_1 _12603_ (.A1(net3627),
    .A2(net380),
    .B1(net358),
    .B2(_02774_),
    .X(_06325_));
 sky130_fd_sc_hd__a21o_1 _12604_ (.A1(_02840_),
    .A2(net378),
    .B1(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__a21oi_4 _12605_ (.A1(net360),
    .A2(_06326_),
    .B1(_06324_),
    .Y(_06327_));
 sky130_fd_sc_hd__o21a_1 _12606_ (.A1(net478),
    .A2(_06327_),
    .B1(_02844_),
    .X(_06328_));
 sky130_fd_sc_hd__nor2_1 _12607_ (.A(net891),
    .B(_06328_),
    .Y(_01164_));
 sky130_fd_sc_hd__mux4_1 _12608_ (.A0(\dpath.RF.R[24][12] ),
    .A1(\dpath.RF.R[25][12] ),
    .A2(\dpath.RF.R[26][12] ),
    .A3(\dpath.RF.R[27][12] ),
    .S0(net823),
    .S1(net803),
    .X(_06329_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(\dpath.RF.R[30][12] ),
    .A1(\dpath.RF.R[31][12] ),
    .S(net824),
    .X(_06330_));
 sky130_fd_sc_hd__mux2_1 _12610_ (.A0(\dpath.RF.R[28][12] ),
    .A1(\dpath.RF.R[29][12] ),
    .S(net831),
    .X(_06331_));
 sky130_fd_sc_hd__a21o_1 _12611_ (.A1(net502),
    .A2(_06331_),
    .B1(net496),
    .X(_06332_));
 sky130_fd_sc_hd__a21o_1 _12612_ (.A1(net803),
    .A2(_06330_),
    .B1(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__o211a_1 _12613_ (.A1(net796),
    .A2(_06329_),
    .B1(_06333_),
    .C1(net794),
    .X(_06334_));
 sky130_fd_sc_hd__mux4_1 _12614_ (.A0(net1506),
    .A1(net2828),
    .A2(net1450),
    .A3(net2698),
    .S0(net823),
    .S1(net803),
    .X(_06335_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(net2760),
    .A1(net2422),
    .S(net824),
    .X(_06336_));
 sky130_fd_sc_hd__mux2_1 _12616_ (.A0(\dpath.RF.R[16][12] ),
    .A1(\dpath.RF.R[17][12] ),
    .S(net831),
    .X(_06337_));
 sky130_fd_sc_hd__a21o_1 _12617_ (.A1(net502),
    .A2(_06337_),
    .B1(net796),
    .X(_06338_));
 sky130_fd_sc_hd__a21o_1 _12618_ (.A1(net803),
    .A2(_06336_),
    .B1(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__o211a_1 _12619_ (.A1(net496),
    .A2(_06335_),
    .B1(_06339_),
    .C1(net491),
    .X(_06340_));
 sky130_fd_sc_hd__or3b_1 _12620_ (.A(_06334_),
    .B(_06340_),
    .C_N(net790),
    .X(_06341_));
 sky130_fd_sc_hd__mux4_1 _12621_ (.A0(\dpath.RF.R[12][12] ),
    .A1(\dpath.RF.R[13][12] ),
    .A2(\dpath.RF.R[14][12] ),
    .A3(\dpath.RF.R[15][12] ),
    .S0(net823),
    .S1(net803),
    .X(_06342_));
 sky130_fd_sc_hd__mux4_1 _12622_ (.A0(\dpath.RF.R[8][12] ),
    .A1(\dpath.RF.R[9][12] ),
    .A2(\dpath.RF.R[10][12] ),
    .A3(\dpath.RF.R[11][12] ),
    .S0(net823),
    .S1(net803),
    .X(_06343_));
 sky130_fd_sc_hd__mux4_1 _12623_ (.A0(\dpath.RF.R[0][12] ),
    .A1(\dpath.RF.R[1][12] ),
    .A2(\dpath.RF.R[2][12] ),
    .A3(\dpath.RF.R[3][12] ),
    .S0(net823),
    .S1(net803),
    .X(_06344_));
 sky130_fd_sc_hd__mux4_1 _12624_ (.A0(\dpath.RF.R[4][12] ),
    .A1(\dpath.RF.R[5][12] ),
    .A2(\dpath.RF.R[6][12] ),
    .A3(\dpath.RF.R[7][12] ),
    .S0(net823),
    .S1(net803),
    .X(_06345_));
 sky130_fd_sc_hd__mux4_1 _12625_ (.A0(_06342_),
    .A1(_06343_),
    .A2(_06345_),
    .A3(_06344_),
    .S0(net496),
    .S1(net491),
    .X(_06346_));
 sky130_fd_sc_hd__or2_1 _12626_ (.A(net790),
    .B(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__and3_1 _12627_ (.A(net364),
    .B(_06341_),
    .C(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__a22o_1 _12628_ (.A1(net694),
    .A2(net380),
    .B1(net358),
    .B2(_02874_),
    .X(_06349_));
 sky130_fd_sc_hd__a21o_1 _12629_ (.A1(_02944_),
    .A2(net378),
    .B1(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__a21oi_4 _12630_ (.A1(net360),
    .A2(_06350_),
    .B1(_06348_),
    .Y(_06351_));
 sky130_fd_sc_hd__o21a_1 _12631_ (.A1(net477),
    .A2(_06351_),
    .B1(net472),
    .X(_06352_));
 sky130_fd_sc_hd__nor2_1 _12632_ (.A(net888),
    .B(_06352_),
    .Y(_01165_));
 sky130_fd_sc_hd__mux4_1 _12633_ (.A0(\dpath.RF.R[24][13] ),
    .A1(\dpath.RF.R[25][13] ),
    .A2(\dpath.RF.R[26][13] ),
    .A3(\dpath.RF.R[27][13] ),
    .S0(net822),
    .S1(net802),
    .X(_06353_));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(\dpath.RF.R[30][13] ),
    .A1(\dpath.RF.R[31][13] ),
    .S(net824),
    .X(_06354_));
 sky130_fd_sc_hd__mux2_1 _12635_ (.A0(\dpath.RF.R[28][13] ),
    .A1(\dpath.RF.R[29][13] ),
    .S(net824),
    .X(_06355_));
 sky130_fd_sc_hd__a21o_1 _12636_ (.A1(net502),
    .A2(_06355_),
    .B1(net496),
    .X(_06356_));
 sky130_fd_sc_hd__a21o_1 _12637_ (.A1(net804),
    .A2(_06354_),
    .B1(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__o211a_1 _12638_ (.A1(net796),
    .A2(_06353_),
    .B1(_06357_),
    .C1(net794),
    .X(_06358_));
 sky130_fd_sc_hd__mux4_1 _12639_ (.A0(\dpath.RF.R[20][13] ),
    .A1(\dpath.RF.R[21][13] ),
    .A2(\dpath.RF.R[22][13] ),
    .A3(\dpath.RF.R[23][13] ),
    .S0(net824),
    .S1(net804),
    .X(_06359_));
 sky130_fd_sc_hd__mux2_1 _12640_ (.A0(\dpath.RF.R[18][13] ),
    .A1(\dpath.RF.R[19][13] ),
    .S(net824),
    .X(_06360_));
 sky130_fd_sc_hd__mux2_1 _12641_ (.A0(\dpath.RF.R[16][13] ),
    .A1(\dpath.RF.R[17][13] ),
    .S(net824),
    .X(_06361_));
 sky130_fd_sc_hd__a21o_1 _12642_ (.A1(net502),
    .A2(_06361_),
    .B1(net796),
    .X(_06362_));
 sky130_fd_sc_hd__a21o_1 _12643_ (.A1(net802),
    .A2(_06360_),
    .B1(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__o211a_1 _12644_ (.A1(net495),
    .A2(_06359_),
    .B1(_06363_),
    .C1(net491),
    .X(_06364_));
 sky130_fd_sc_hd__or3b_1 _12645_ (.A(_06358_),
    .B(_06364_),
    .C_N(net790),
    .X(_06365_));
 sky130_fd_sc_hd__mux4_1 _12646_ (.A0(\dpath.RF.R[12][13] ),
    .A1(\dpath.RF.R[13][13] ),
    .A2(\dpath.RF.R[14][13] ),
    .A3(\dpath.RF.R[15][13] ),
    .S0(net824),
    .S1(net802),
    .X(_06366_));
 sky130_fd_sc_hd__mux4_1 _12647_ (.A0(\dpath.RF.R[8][13] ),
    .A1(\dpath.RF.R[9][13] ),
    .A2(\dpath.RF.R[10][13] ),
    .A3(\dpath.RF.R[11][13] ),
    .S0(net824),
    .S1(net804),
    .X(_06367_));
 sky130_fd_sc_hd__mux4_1 _12648_ (.A0(\dpath.RF.R[0][13] ),
    .A1(\dpath.RF.R[1][13] ),
    .A2(\dpath.RF.R[2][13] ),
    .A3(\dpath.RF.R[3][13] ),
    .S0(net822),
    .S1(net802),
    .X(_06368_));
 sky130_fd_sc_hd__mux4_1 _12649_ (.A0(\dpath.RF.R[4][13] ),
    .A1(\dpath.RF.R[5][13] ),
    .A2(\dpath.RF.R[6][13] ),
    .A3(\dpath.RF.R[7][13] ),
    .S0(net822),
    .S1(net802),
    .X(_06369_));
 sky130_fd_sc_hd__mux4_1 _12650_ (.A0(_06366_),
    .A1(_06367_),
    .A2(_06369_),
    .A3(_06368_),
    .S0(net496),
    .S1(net491),
    .X(_06370_));
 sky130_fd_sc_hd__or2_1 _12651_ (.A(net790),
    .B(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__and3_1 _12652_ (.A(net364),
    .B(_06365_),
    .C(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__a22o_1 _12653_ (.A1(net693),
    .A2(net380),
    .B1(net358),
    .B2(_02977_),
    .X(_06373_));
 sky130_fd_sc_hd__a21o_1 _12654_ (.A1(_03052_),
    .A2(net378),
    .B1(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__a21oi_4 _12655_ (.A1(net360),
    .A2(_06374_),
    .B1(_06372_),
    .Y(_06375_));
 sky130_fd_sc_hd__o21a_1 _12656_ (.A1(net477),
    .A2(_06375_),
    .B1(net472),
    .X(_06376_));
 sky130_fd_sc_hd__nor2_1 _12657_ (.A(net888),
    .B(_06376_),
    .Y(_01166_));
 sky130_fd_sc_hd__mux4_1 _12658_ (.A0(net1804),
    .A1(net1548),
    .A2(net1910),
    .A3(net2192),
    .S0(net826),
    .S1(net806),
    .X(_06377_));
 sky130_fd_sc_hd__mux2_1 _12659_ (.A0(net2290),
    .A1(net2976),
    .S(net836),
    .X(_06378_));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(\dpath.RF.R[28][14] ),
    .A1(\dpath.RF.R[29][14] ),
    .S(net836),
    .X(_06379_));
 sky130_fd_sc_hd__a21o_1 _12661_ (.A1(net503),
    .A2(_06379_),
    .B1(net497),
    .X(_06380_));
 sky130_fd_sc_hd__a21o_1 _12662_ (.A1(net806),
    .A2(_06378_),
    .B1(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__o211a_1 _12663_ (.A1(net797),
    .A2(_06377_),
    .B1(_06381_),
    .C1(net794),
    .X(_06382_));
 sky130_fd_sc_hd__mux4_1 _12664_ (.A0(net1694),
    .A1(net3693),
    .A2(net1596),
    .A3(net2450),
    .S0(net826),
    .S1(net806),
    .X(_06383_));
 sky130_fd_sc_hd__mux2_1 _12665_ (.A0(net2728),
    .A1(net2706),
    .S(net826),
    .X(_06384_));
 sky130_fd_sc_hd__mux2_1 _12666_ (.A0(\dpath.RF.R[16][14] ),
    .A1(\dpath.RF.R[17][14] ),
    .S(net836),
    .X(_06385_));
 sky130_fd_sc_hd__a21o_1 _12667_ (.A1(net503),
    .A2(_06385_),
    .B1(net797),
    .X(_06386_));
 sky130_fd_sc_hd__a21o_1 _12668_ (.A1(net806),
    .A2(_06384_),
    .B1(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__o211a_1 _12669_ (.A1(net497),
    .A2(_06383_),
    .B1(_06387_),
    .C1(net492),
    .X(_06388_));
 sky130_fd_sc_hd__or3b_1 _12670_ (.A(_06382_),
    .B(_06388_),
    .C_N(net791),
    .X(_06389_));
 sky130_fd_sc_hd__mux4_1 _12671_ (.A0(\dpath.RF.R[12][14] ),
    .A1(\dpath.RF.R[13][14] ),
    .A2(\dpath.RF.R[14][14] ),
    .A3(\dpath.RF.R[15][14] ),
    .S0(net831),
    .S1(net810),
    .X(_06390_));
 sky130_fd_sc_hd__mux4_1 _12672_ (.A0(\dpath.RF.R[8][14] ),
    .A1(\dpath.RF.R[9][14] ),
    .A2(\dpath.RF.R[10][14] ),
    .A3(\dpath.RF.R[11][14] ),
    .S0(net824),
    .S1(net803),
    .X(_06391_));
 sky130_fd_sc_hd__mux4_1 _12673_ (.A0(\dpath.RF.R[0][14] ),
    .A1(\dpath.RF.R[1][14] ),
    .A2(\dpath.RF.R[2][14] ),
    .A3(\dpath.RF.R[3][14] ),
    .S0(net823),
    .S1(net803),
    .X(_06392_));
 sky130_fd_sc_hd__mux4_1 _12674_ (.A0(\dpath.RF.R[4][14] ),
    .A1(\dpath.RF.R[5][14] ),
    .A2(\dpath.RF.R[6][14] ),
    .A3(\dpath.RF.R[7][14] ),
    .S0(net823),
    .S1(net803),
    .X(_06393_));
 sky130_fd_sc_hd__mux4_1 _12675_ (.A0(_06390_),
    .A1(_06391_),
    .A2(_06393_),
    .A3(_06392_),
    .S0(net496),
    .S1(net491),
    .X(_06394_));
 sky130_fd_sc_hd__or2_1 _12676_ (.A(net790),
    .B(_06394_),
    .X(_06395_));
 sky130_fd_sc_hd__and3_1 _12677_ (.A(net364),
    .B(_06389_),
    .C(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__a22o_1 _12678_ (.A1(net690),
    .A2(net379),
    .B1(net357),
    .B2(_03087_),
    .X(_06397_));
 sky130_fd_sc_hd__a21o_1 _12679_ (.A1(_03166_),
    .A2(net378),
    .B1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a21oi_4 _12680_ (.A1(net359),
    .A2(_06398_),
    .B1(_06396_),
    .Y(_06399_));
 sky130_fd_sc_hd__o21a_1 _12681_ (.A1(net477),
    .A2(_06399_),
    .B1(net472),
    .X(_06400_));
 sky130_fd_sc_hd__nor2_1 _12682_ (.A(net888),
    .B(_06400_),
    .Y(_01167_));
 sky130_fd_sc_hd__mux4_1 _12683_ (.A0(\dpath.RF.R[24][15] ),
    .A1(\dpath.RF.R[25][15] ),
    .A2(\dpath.RF.R[26][15] ),
    .A3(\dpath.RF.R[27][15] ),
    .S0(net822),
    .S1(net802),
    .X(_06401_));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(\dpath.RF.R[30][15] ),
    .A1(\dpath.RF.R[31][15] ),
    .S(net831),
    .X(_06402_));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(\dpath.RF.R[28][15] ),
    .A1(\dpath.RF.R[29][15] ),
    .S(net831),
    .X(_06403_));
 sky130_fd_sc_hd__a21o_1 _12686_ (.A1(net503),
    .A2(_06403_),
    .B1(net496),
    .X(_06404_));
 sky130_fd_sc_hd__a21o_1 _12687_ (.A1(net804),
    .A2(_06402_),
    .B1(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__o211a_1 _12688_ (.A1(net797),
    .A2(_06401_),
    .B1(_06405_),
    .C1(net794),
    .X(_06406_));
 sky130_fd_sc_hd__mux4_1 _12689_ (.A0(net1652),
    .A1(\dpath.RF.R[21][15] ),
    .A2(\dpath.RF.R[22][15] ),
    .A3(\dpath.RF.R[23][15] ),
    .S0(net822),
    .S1(net804),
    .X(_06407_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(net1642),
    .A1(\dpath.RF.R[19][15] ),
    .S(net830),
    .X(_06408_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(\dpath.RF.R[16][15] ),
    .A1(\dpath.RF.R[17][15] ),
    .S(net830),
    .X(_06409_));
 sky130_fd_sc_hd__a21o_1 _12692_ (.A1(net503),
    .A2(_06409_),
    .B1(net797),
    .X(_06410_));
 sky130_fd_sc_hd__a21o_1 _12693_ (.A1(net802),
    .A2(_06408_),
    .B1(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__o211a_1 _12694_ (.A1(net496),
    .A2(_06407_),
    .B1(_06411_),
    .C1(net492),
    .X(_06412_));
 sky130_fd_sc_hd__or3b_1 _12695_ (.A(_06406_),
    .B(_06412_),
    .C_N(net792),
    .X(_06413_));
 sky130_fd_sc_hd__mux4_1 _12696_ (.A0(\dpath.RF.R[12][15] ),
    .A1(\dpath.RF.R[13][15] ),
    .A2(\dpath.RF.R[14][15] ),
    .A3(\dpath.RF.R[15][15] ),
    .S0(net830),
    .S1(net809),
    .X(_06414_));
 sky130_fd_sc_hd__mux4_1 _12697_ (.A0(\dpath.RF.R[8][15] ),
    .A1(\dpath.RF.R[9][15] ),
    .A2(\dpath.RF.R[10][15] ),
    .A3(\dpath.RF.R[11][15] ),
    .S0(net822),
    .S1(net802),
    .X(_06415_));
 sky130_fd_sc_hd__mux4_1 _12698_ (.A0(\dpath.RF.R[0][15] ),
    .A1(\dpath.RF.R[1][15] ),
    .A2(\dpath.RF.R[2][15] ),
    .A3(\dpath.RF.R[3][15] ),
    .S0(net822),
    .S1(net802),
    .X(_06416_));
 sky130_fd_sc_hd__mux4_1 _12699_ (.A0(\dpath.RF.R[4][15] ),
    .A1(\dpath.RF.R[5][15] ),
    .A2(\dpath.RF.R[6][15] ),
    .A3(\dpath.RF.R[7][15] ),
    .S0(net822),
    .S1(net802),
    .X(_06417_));
 sky130_fd_sc_hd__mux4_1 _12700_ (.A0(_06414_),
    .A1(_06415_),
    .A2(_06417_),
    .A3(_06416_),
    .S0(net496),
    .S1(net492),
    .X(_06418_));
 sky130_fd_sc_hd__or2_1 _12701_ (.A(net792),
    .B(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__and3_1 _12702_ (.A(net363),
    .B(_06413_),
    .C(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__a22o_1 _12703_ (.A1(net688),
    .A2(net379),
    .B1(net357),
    .B2(_03198_),
    .X(_06421_));
 sky130_fd_sc_hd__a21o_1 _12704_ (.A1(_03282_),
    .A2(net377),
    .B1(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__a21oi_4 _12705_ (.A1(net359),
    .A2(_06422_),
    .B1(_06420_),
    .Y(_06423_));
 sky130_fd_sc_hd__o21a_1 _12706_ (.A1(net477),
    .A2(_06423_),
    .B1(net472),
    .X(_06424_));
 sky130_fd_sc_hd__nor2_1 _12707_ (.A(net888),
    .B(_06424_),
    .Y(_01168_));
 sky130_fd_sc_hd__mux4_1 _12708_ (.A0(net1300),
    .A1(\dpath.RF.R[25][16] ),
    .A2(\dpath.RF.R[26][16] ),
    .A3(\dpath.RF.R[27][16] ),
    .S0(net830),
    .S1(net809),
    .X(_06425_));
 sky130_fd_sc_hd__mux2_1 _12709_ (.A0(net1290),
    .A1(\dpath.RF.R[31][16] ),
    .S(net832),
    .X(_06426_));
 sky130_fd_sc_hd__mux2_1 _12710_ (.A0(\dpath.RF.R[28][16] ),
    .A1(\dpath.RF.R[29][16] ),
    .S(net830),
    .X(_06427_));
 sky130_fd_sc_hd__a21o_1 _12711_ (.A1(net504),
    .A2(_06427_),
    .B1(net498),
    .X(_06428_));
 sky130_fd_sc_hd__a21o_1 _12712_ (.A1(net809),
    .A2(_06426_),
    .B1(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__o211a_1 _12713_ (.A1(net798),
    .A2(_06425_),
    .B1(_06429_),
    .C1(net795),
    .X(_06430_));
 sky130_fd_sc_hd__mux4_1 _12714_ (.A0(net3705),
    .A1(\dpath.RF.R[21][16] ),
    .A2(\dpath.RF.R[22][16] ),
    .A3(net2518),
    .S0(net830),
    .S1(net809),
    .X(_06431_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(\dpath.RF.R[18][16] ),
    .A1(\dpath.RF.R[19][16] ),
    .S(net830),
    .X(_06432_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(\dpath.RF.R[16][16] ),
    .A1(\dpath.RF.R[17][16] ),
    .S(net832),
    .X(_06433_));
 sky130_fd_sc_hd__a21o_1 _12717_ (.A1(net504),
    .A2(_06433_),
    .B1(net798),
    .X(_06434_));
 sky130_fd_sc_hd__a21o_1 _12718_ (.A1(net809),
    .A2(_06432_),
    .B1(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__o211a_1 _12719_ (.A1(net498),
    .A2(_06431_),
    .B1(_06435_),
    .C1(net493),
    .X(_06436_));
 sky130_fd_sc_hd__or3b_1 _12720_ (.A(_06430_),
    .B(_06436_),
    .C_N(net793),
    .X(_06437_));
 sky130_fd_sc_hd__mux4_1 _12721_ (.A0(\dpath.RF.R[12][16] ),
    .A1(\dpath.RF.R[13][16] ),
    .A2(\dpath.RF.R[14][16] ),
    .A3(\dpath.RF.R[15][16] ),
    .S0(net832),
    .S1(net809),
    .X(_06438_));
 sky130_fd_sc_hd__mux4_1 _12722_ (.A0(\dpath.RF.R[8][16] ),
    .A1(\dpath.RF.R[9][16] ),
    .A2(\dpath.RF.R[10][16] ),
    .A3(\dpath.RF.R[11][16] ),
    .S0(net830),
    .S1(net809),
    .X(_06439_));
 sky130_fd_sc_hd__mux4_1 _12723_ (.A0(\dpath.RF.R[0][16] ),
    .A1(\dpath.RF.R[1][16] ),
    .A2(\dpath.RF.R[2][16] ),
    .A3(\dpath.RF.R[3][16] ),
    .S0(net832),
    .S1(net809),
    .X(_06440_));
 sky130_fd_sc_hd__mux4_1 _12724_ (.A0(\dpath.RF.R[4][16] ),
    .A1(\dpath.RF.R[5][16] ),
    .A2(\dpath.RF.R[6][16] ),
    .A3(\dpath.RF.R[7][16] ),
    .S0(net832),
    .S1(net810),
    .X(_06441_));
 sky130_fd_sc_hd__mux4_1 _12725_ (.A0(_06438_),
    .A1(_06439_),
    .A2(_06441_),
    .A3(_06440_),
    .S0(net498),
    .S1(net493),
    .X(_06442_));
 sky130_fd_sc_hd__or2_1 _12726_ (.A(net792),
    .B(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__and3_1 _12727_ (.A(net363),
    .B(_06437_),
    .C(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__a22o_1 _12728_ (.A1(net686),
    .A2(net379),
    .B1(net357),
    .B2(_03317_),
    .X(_06445_));
 sky130_fd_sc_hd__a21o_1 _12729_ (.A1(_03411_),
    .A2(net377),
    .B1(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__a21oi_4 _12730_ (.A1(net359),
    .A2(_06446_),
    .B1(_06444_),
    .Y(_06447_));
 sky130_fd_sc_hd__o21a_1 _12731_ (.A1(net477),
    .A2(_06447_),
    .B1(net472),
    .X(_06448_));
 sky130_fd_sc_hd__nor2_1 _12732_ (.A(net885),
    .B(_06448_),
    .Y(_01169_));
 sky130_fd_sc_hd__mux4_1 _12733_ (.A0(\dpath.RF.R[24][17] ),
    .A1(\dpath.RF.R[25][17] ),
    .A2(\dpath.RF.R[26][17] ),
    .A3(\dpath.RF.R[27][17] ),
    .S0(net830),
    .S1(net809),
    .X(_06449_));
 sky130_fd_sc_hd__mux2_1 _12734_ (.A0(\dpath.RF.R[30][17] ),
    .A1(\dpath.RF.R[31][17] ),
    .S(net831),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_1 _12735_ (.A0(\dpath.RF.R[28][17] ),
    .A1(\dpath.RF.R[29][17] ),
    .S(net831),
    .X(_06451_));
 sky130_fd_sc_hd__a21o_1 _12736_ (.A1(net504),
    .A2(_06451_),
    .B1(net498),
    .X(_06452_));
 sky130_fd_sc_hd__a21o_1 _12737_ (.A1(net809),
    .A2(_06450_),
    .B1(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__o211a_1 _12738_ (.A1(net798),
    .A2(_06449_),
    .B1(_06453_),
    .C1(net795),
    .X(_06454_));
 sky130_fd_sc_hd__mux4_1 _12739_ (.A0(\dpath.RF.R[20][17] ),
    .A1(net2098),
    .A2(net3700),
    .A3(net1768),
    .S0(net830),
    .S1(net809),
    .X(_06455_));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(net1872),
    .A1(\dpath.RF.R[19][17] ),
    .S(net830),
    .X(_06456_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(\dpath.RF.R[16][17] ),
    .A1(\dpath.RF.R[17][17] ),
    .S(net830),
    .X(_06457_));
 sky130_fd_sc_hd__a21o_1 _12742_ (.A1(net504),
    .A2(_06457_),
    .B1(net798),
    .X(_06458_));
 sky130_fd_sc_hd__a21o_1 _12743_ (.A1(net809),
    .A2(_06456_),
    .B1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__o211a_1 _12744_ (.A1(net498),
    .A2(net3701),
    .B1(_06459_),
    .C1(net493),
    .X(_06460_));
 sky130_fd_sc_hd__or3b_1 _12745_ (.A(_06454_),
    .B(net3702),
    .C_N(net792),
    .X(_06461_));
 sky130_fd_sc_hd__mux4_1 _12746_ (.A0(\dpath.RF.R[12][17] ),
    .A1(\dpath.RF.R[13][17] ),
    .A2(\dpath.RF.R[14][17] ),
    .A3(\dpath.RF.R[15][17] ),
    .S0(net830),
    .S1(net809),
    .X(_06462_));
 sky130_fd_sc_hd__mux4_1 _12747_ (.A0(\dpath.RF.R[8][17] ),
    .A1(\dpath.RF.R[9][17] ),
    .A2(\dpath.RF.R[10][17] ),
    .A3(\dpath.RF.R[11][17] ),
    .S0(net830),
    .S1(net809),
    .X(_06463_));
 sky130_fd_sc_hd__mux4_1 _12748_ (.A0(\dpath.RF.R[0][17] ),
    .A1(\dpath.RF.R[1][17] ),
    .A2(\dpath.RF.R[2][17] ),
    .A3(\dpath.RF.R[3][17] ),
    .S0(net830),
    .S1(net809),
    .X(_06464_));
 sky130_fd_sc_hd__mux4_1 _12749_ (.A0(\dpath.RF.R[4][17] ),
    .A1(\dpath.RF.R[5][17] ),
    .A2(\dpath.RF.R[6][17] ),
    .A3(\dpath.RF.R[7][17] ),
    .S0(net830),
    .S1(net809),
    .X(_06465_));
 sky130_fd_sc_hd__mux4_1 _12750_ (.A0(_06462_),
    .A1(_06463_),
    .A2(_06465_),
    .A3(_06464_),
    .S0(net498),
    .S1(net493),
    .X(_06466_));
 sky130_fd_sc_hd__or2_1 _12751_ (.A(net792),
    .B(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__and3_1 _12752_ (.A(net363),
    .B(_06461_),
    .C(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__a22o_1 _12753_ (.A1(net684),
    .A2(net379),
    .B1(net357),
    .B2(_03445_),
    .X(_06469_));
 sky130_fd_sc_hd__a21o_1 _12754_ (.A1(_03543_),
    .A2(net377),
    .B1(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__a21oi_4 _12755_ (.A1(net359),
    .A2(_06470_),
    .B1(_06468_),
    .Y(_06471_));
 sky130_fd_sc_hd__o21a_1 _12756_ (.A1(net477),
    .A2(_06471_),
    .B1(net472),
    .X(_06472_));
 sky130_fd_sc_hd__nor2_1 _12757_ (.A(net886),
    .B(_06472_),
    .Y(_01170_));
 sky130_fd_sc_hd__mux4_1 _12758_ (.A0(\dpath.RF.R[24][18] ),
    .A1(\dpath.RF.R[25][18] ),
    .A2(\dpath.RF.R[26][18] ),
    .A3(\dpath.RF.R[27][18] ),
    .S0(net831),
    .S1(net810),
    .X(_06473_));
 sky130_fd_sc_hd__mux2_1 _12759_ (.A0(\dpath.RF.R[30][18] ),
    .A1(\dpath.RF.R[31][18] ),
    .S(net834),
    .X(_06474_));
 sky130_fd_sc_hd__mux2_1 _12760_ (.A0(\dpath.RF.R[28][18] ),
    .A1(\dpath.RF.R[29][18] ),
    .S(net834),
    .X(_06475_));
 sky130_fd_sc_hd__a21o_1 _12761_ (.A1(net504),
    .A2(_06475_),
    .B1(net498),
    .X(_06476_));
 sky130_fd_sc_hd__a21o_1 _12762_ (.A1(net812),
    .A2(_06474_),
    .B1(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__o211a_1 _12763_ (.A1(net798),
    .A2(_06473_),
    .B1(_06477_),
    .C1(net795),
    .X(_06478_));
 sky130_fd_sc_hd__mux4_1 _12764_ (.A0(net1568),
    .A1(\dpath.RF.R[21][18] ),
    .A2(\dpath.RF.R[22][18] ),
    .A3(\dpath.RF.R[23][18] ),
    .S0(net833),
    .S1(net811),
    .X(_06479_));
 sky130_fd_sc_hd__mux2_1 _12765_ (.A0(net1478),
    .A1(\dpath.RF.R[19][18] ),
    .S(net833),
    .X(_06480_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(\dpath.RF.R[16][18] ),
    .A1(\dpath.RF.R[17][18] ),
    .S(net833),
    .X(_06481_));
 sky130_fd_sc_hd__a21o_1 _12767_ (.A1(net504),
    .A2(_06481_),
    .B1(net798),
    .X(_06482_));
 sky130_fd_sc_hd__a21o_1 _12768_ (.A1(net811),
    .A2(_06480_),
    .B1(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__o211a_1 _12769_ (.A1(net499),
    .A2(_06479_),
    .B1(_06483_),
    .C1(net493),
    .X(_06484_));
 sky130_fd_sc_hd__or3b_1 _12770_ (.A(_06478_),
    .B(_06484_),
    .C_N(net792),
    .X(_06485_));
 sky130_fd_sc_hd__mux4_1 _12771_ (.A0(\dpath.RF.R[12][18] ),
    .A1(\dpath.RF.R[13][18] ),
    .A2(\dpath.RF.R[14][18] ),
    .A3(\dpath.RF.R[15][18] ),
    .S0(net833),
    .S1(net811),
    .X(_06486_));
 sky130_fd_sc_hd__mux4_1 _12772_ (.A0(\dpath.RF.R[8][18] ),
    .A1(\dpath.RF.R[9][18] ),
    .A2(\dpath.RF.R[10][18] ),
    .A3(\dpath.RF.R[11][18] ),
    .S0(net833),
    .S1(net811),
    .X(_06487_));
 sky130_fd_sc_hd__mux4_1 _12773_ (.A0(\dpath.RF.R[0][18] ),
    .A1(\dpath.RF.R[1][18] ),
    .A2(\dpath.RF.R[2][18] ),
    .A3(\dpath.RF.R[3][18] ),
    .S0(net833),
    .S1(net811),
    .X(_06488_));
 sky130_fd_sc_hd__mux4_1 _12774_ (.A0(\dpath.RF.R[4][18] ),
    .A1(\dpath.RF.R[5][18] ),
    .A2(\dpath.RF.R[6][18] ),
    .A3(\dpath.RF.R[7][18] ),
    .S0(net833),
    .S1(net811),
    .X(_06489_));
 sky130_fd_sc_hd__mux4_1 _12775_ (.A0(_06486_),
    .A1(_06487_),
    .A2(_06489_),
    .A3(_06488_),
    .S0(net498),
    .S1(net493),
    .X(_06490_));
 sky130_fd_sc_hd__or2_1 _12776_ (.A(net792),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__and3_1 _12777_ (.A(net363),
    .B(_06485_),
    .C(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__a22o_1 _12778_ (.A1(net683),
    .A2(net379),
    .B1(net357),
    .B2(_03578_),
    .X(_06493_));
 sky130_fd_sc_hd__a21o_1 _12779_ (.A1(_03684_),
    .A2(net377),
    .B1(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__a21oi_4 _12780_ (.A1(net359),
    .A2(_06494_),
    .B1(_06492_),
    .Y(_06495_));
 sky130_fd_sc_hd__o21a_1 _12781_ (.A1(net477),
    .A2(_06495_),
    .B1(net472),
    .X(_06496_));
 sky130_fd_sc_hd__nor2_1 _12782_ (.A(net885),
    .B(_06496_),
    .Y(_01171_));
 sky130_fd_sc_hd__mux4_1 _12783_ (.A0(\dpath.RF.R[24][19] ),
    .A1(\dpath.RF.R[25][19] ),
    .A2(\dpath.RF.R[26][19] ),
    .A3(\dpath.RF.R[27][19] ),
    .S0(net831),
    .S1(net810),
    .X(_06497_));
 sky130_fd_sc_hd__mux2_1 _12784_ (.A0(net1406),
    .A1(\dpath.RF.R[31][19] ),
    .S(net832),
    .X(_06498_));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(\dpath.RF.R[28][19] ),
    .A1(\dpath.RF.R[29][19] ),
    .S(net832),
    .X(_06499_));
 sky130_fd_sc_hd__a21o_1 _12786_ (.A1(net504),
    .A2(_06499_),
    .B1(net498),
    .X(_06500_));
 sky130_fd_sc_hd__a21o_1 _12787_ (.A1(net810),
    .A2(_06498_),
    .B1(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__o211a_1 _12788_ (.A1(net798),
    .A2(_06497_),
    .B1(_06501_),
    .C1(net795),
    .X(_06502_));
 sky130_fd_sc_hd__mux4_1 _12789_ (.A0(\dpath.RF.R[20][19] ),
    .A1(\dpath.RF.R[21][19] ),
    .A2(\dpath.RF.R[22][19] ),
    .A3(\dpath.RF.R[23][19] ),
    .S0(net831),
    .S1(net810),
    .X(_06503_));
 sky130_fd_sc_hd__mux2_1 _12790_ (.A0(\dpath.RF.R[18][19] ),
    .A1(\dpath.RF.R[19][19] ),
    .S(net832),
    .X(_06504_));
 sky130_fd_sc_hd__mux2_1 _12791_ (.A0(\dpath.RF.R[16][19] ),
    .A1(\dpath.RF.R[17][19] ),
    .S(net832),
    .X(_06505_));
 sky130_fd_sc_hd__a21o_1 _12792_ (.A1(net504),
    .A2(_06505_),
    .B1(net798),
    .X(_06506_));
 sky130_fd_sc_hd__a21o_1 _12793_ (.A1(net810),
    .A2(_06504_),
    .B1(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__o211a_1 _12794_ (.A1(net498),
    .A2(_06503_),
    .B1(_06507_),
    .C1(net493),
    .X(_06508_));
 sky130_fd_sc_hd__or3b_1 _12795_ (.A(_06502_),
    .B(_06508_),
    .C_N(net792),
    .X(_06509_));
 sky130_fd_sc_hd__mux4_1 _12796_ (.A0(\dpath.RF.R[12][19] ),
    .A1(\dpath.RF.R[13][19] ),
    .A2(\dpath.RF.R[14][19] ),
    .A3(\dpath.RF.R[15][19] ),
    .S0(net832),
    .S1(net810),
    .X(_06510_));
 sky130_fd_sc_hd__mux4_1 _12797_ (.A0(\dpath.RF.R[8][19] ),
    .A1(\dpath.RF.R[9][19] ),
    .A2(\dpath.RF.R[10][19] ),
    .A3(\dpath.RF.R[11][19] ),
    .S0(net831),
    .S1(net810),
    .X(_06511_));
 sky130_fd_sc_hd__mux4_1 _12798_ (.A0(\dpath.RF.R[0][19] ),
    .A1(\dpath.RF.R[1][19] ),
    .A2(\dpath.RF.R[2][19] ),
    .A3(\dpath.RF.R[3][19] ),
    .S0(net831),
    .S1(net810),
    .X(_06512_));
 sky130_fd_sc_hd__mux4_1 _12799_ (.A0(\dpath.RF.R[4][19] ),
    .A1(\dpath.RF.R[5][19] ),
    .A2(\dpath.RF.R[6][19] ),
    .A3(\dpath.RF.R[7][19] ),
    .S0(net831),
    .S1(net810),
    .X(_06513_));
 sky130_fd_sc_hd__mux4_1 _12800_ (.A0(_06510_),
    .A1(_06511_),
    .A2(_06513_),
    .A3(_06512_),
    .S0(net498),
    .S1(net493),
    .X(_06514_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(net792),
    .B(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__and3_1 _12802_ (.A(net363),
    .B(_06509_),
    .C(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__a22o_1 _12803_ (.A1(net680),
    .A2(net379),
    .B1(net357),
    .B2(_03719_),
    .X(_06517_));
 sky130_fd_sc_hd__a21o_1 _12804_ (.A1(_03820_),
    .A2(net377),
    .B1(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__a21oi_4 _12805_ (.A1(net359),
    .A2(_06518_),
    .B1(_06516_),
    .Y(_06519_));
 sky130_fd_sc_hd__o21a_1 _12806_ (.A1(net477),
    .A2(_06519_),
    .B1(net472),
    .X(_06520_));
 sky130_fd_sc_hd__nor2_1 _12807_ (.A(net886),
    .B(_06520_),
    .Y(_01172_));
 sky130_fd_sc_hd__mux4_1 _12808_ (.A0(net2614),
    .A1(\dpath.RF.R[25][20] ),
    .A2(\dpath.RF.R[26][20] ),
    .A3(net2068),
    .S0(net833),
    .S1(net811),
    .X(_06521_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(net1810),
    .A1(\dpath.RF.R[31][20] ),
    .S(net833),
    .X(_06522_));
 sky130_fd_sc_hd__mux2_1 _12810_ (.A0(\dpath.RF.R[28][20] ),
    .A1(\dpath.RF.R[29][20] ),
    .S(net833),
    .X(_06523_));
 sky130_fd_sc_hd__a21o_1 _12811_ (.A1(net504),
    .A2(_06523_),
    .B1(net498),
    .X(_06524_));
 sky130_fd_sc_hd__a21o_1 _12812_ (.A1(net811),
    .A2(_06522_),
    .B1(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__o211a_1 _12813_ (.A1(net798),
    .A2(_06521_),
    .B1(_06525_),
    .C1(net795),
    .X(_06526_));
 sky130_fd_sc_hd__mux4_1 _12814_ (.A0(net1700),
    .A1(\dpath.RF.R[21][20] ),
    .A2(net1410),
    .A3(net2658),
    .S0(net833),
    .S1(net811),
    .X(_06527_));
 sky130_fd_sc_hd__mux2_1 _12815_ (.A0(net1538),
    .A1(net1836),
    .S(net835),
    .X(_06528_));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(\dpath.RF.R[16][20] ),
    .A1(\dpath.RF.R[17][20] ),
    .S(net833),
    .X(_06529_));
 sky130_fd_sc_hd__a21o_1 _12817_ (.A1(net504),
    .A2(_06529_),
    .B1(net798),
    .X(_06530_));
 sky130_fd_sc_hd__a21o_1 _12818_ (.A1(net811),
    .A2(_06528_),
    .B1(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__o211a_1 _12819_ (.A1(net498),
    .A2(_06527_),
    .B1(_06531_),
    .C1(net493),
    .X(_06532_));
 sky130_fd_sc_hd__or3b_1 _12820_ (.A(_06526_),
    .B(_06532_),
    .C_N(net792),
    .X(_06533_));
 sky130_fd_sc_hd__mux4_1 _12821_ (.A0(\dpath.RF.R[12][20] ),
    .A1(\dpath.RF.R[13][20] ),
    .A2(\dpath.RF.R[14][20] ),
    .A3(\dpath.RF.R[15][20] ),
    .S0(net835),
    .S1(net813),
    .X(_06534_));
 sky130_fd_sc_hd__mux4_1 _12822_ (.A0(\dpath.RF.R[8][20] ),
    .A1(\dpath.RF.R[9][20] ),
    .A2(\dpath.RF.R[10][20] ),
    .A3(\dpath.RF.R[11][20] ),
    .S0(net835),
    .S1(net811),
    .X(_06535_));
 sky130_fd_sc_hd__mux4_1 _12823_ (.A0(\dpath.RF.R[0][20] ),
    .A1(\dpath.RF.R[1][20] ),
    .A2(\dpath.RF.R[2][20] ),
    .A3(\dpath.RF.R[3][20] ),
    .S0(net833),
    .S1(net811),
    .X(_06536_));
 sky130_fd_sc_hd__mux4_1 _12824_ (.A0(\dpath.RF.R[4][20] ),
    .A1(\dpath.RF.R[5][20] ),
    .A2(\dpath.RF.R[6][20] ),
    .A3(\dpath.RF.R[7][20] ),
    .S0(net835),
    .S1(net813),
    .X(_06537_));
 sky130_fd_sc_hd__mux4_1 _12825_ (.A0(_06534_),
    .A1(_06535_),
    .A2(_06537_),
    .A3(_06536_),
    .S0(net498),
    .S1(net493),
    .X(_06538_));
 sky130_fd_sc_hd__or2_1 _12826_ (.A(net792),
    .B(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__and3_1 _12827_ (.A(net363),
    .B(_06533_),
    .C(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__a22o_1 _12828_ (.A1(net679),
    .A2(net379),
    .B1(net357),
    .B2(_03851_),
    .X(_06541_));
 sky130_fd_sc_hd__a21o_1 _12829_ (.A1(_03968_),
    .A2(net377),
    .B1(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__a21oi_4 _12830_ (.A1(net359),
    .A2(_06542_),
    .B1(_06540_),
    .Y(_06543_));
 sky130_fd_sc_hd__o21a_1 _12831_ (.A1(net477),
    .A2(_06543_),
    .B1(net472),
    .X(_06544_));
 sky130_fd_sc_hd__nor2_1 _12832_ (.A(net885),
    .B(_06544_),
    .Y(_01173_));
 sky130_fd_sc_hd__mux4_1 _12833_ (.A0(net2708),
    .A1(\dpath.RF.R[25][21] ),
    .A2(net3706),
    .A3(net2334),
    .S0(net834),
    .S1(net812),
    .X(_06545_));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(\dpath.RF.R[30][21] ),
    .A1(\dpath.RF.R[31][21] ),
    .S(net834),
    .X(_06546_));
 sky130_fd_sc_hd__mux2_1 _12835_ (.A0(\dpath.RF.R[28][21] ),
    .A1(\dpath.RF.R[29][21] ),
    .S(net835),
    .X(_06547_));
 sky130_fd_sc_hd__a21o_1 _12836_ (.A1(net504),
    .A2(_06547_),
    .B1(net498),
    .X(_06548_));
 sky130_fd_sc_hd__a21o_1 _12837_ (.A1(net813),
    .A2(_06546_),
    .B1(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__o211a_1 _12838_ (.A1(net798),
    .A2(net3707),
    .B1(_06549_),
    .C1(net795),
    .X(_06550_));
 sky130_fd_sc_hd__mux4_1 _12839_ (.A0(net1874),
    .A1(\dpath.RF.R[21][21] ),
    .A2(net1284),
    .A3(net2672),
    .S0(net834),
    .S1(net812),
    .X(_06551_));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(net2022),
    .A1(\dpath.RF.R[19][21] ),
    .S(net833),
    .X(_06552_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(\dpath.RF.R[16][21] ),
    .A1(\dpath.RF.R[17][21] ),
    .S(net833),
    .X(_06553_));
 sky130_fd_sc_hd__a21o_1 _12842_ (.A1(net504),
    .A2(_06553_),
    .B1(net798),
    .X(_06554_));
 sky130_fd_sc_hd__a21o_1 _12843_ (.A1(net813),
    .A2(_06552_),
    .B1(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__o211a_1 _12844_ (.A1(net498),
    .A2(_06551_),
    .B1(_06555_),
    .C1(net493),
    .X(_06556_));
 sky130_fd_sc_hd__or3b_1 _12845_ (.A(_06550_),
    .B(_06556_),
    .C_N(net792),
    .X(_06557_));
 sky130_fd_sc_hd__mux4_1 _12846_ (.A0(\dpath.RF.R[12][21] ),
    .A1(\dpath.RF.R[13][21] ),
    .A2(\dpath.RF.R[14][21] ),
    .A3(\dpath.RF.R[15][21] ),
    .S0(net835),
    .S1(net812),
    .X(_06558_));
 sky130_fd_sc_hd__mux4_1 _12847_ (.A0(\dpath.RF.R[8][21] ),
    .A1(\dpath.RF.R[9][21] ),
    .A2(\dpath.RF.R[10][21] ),
    .A3(\dpath.RF.R[11][21] ),
    .S0(net833),
    .S1(net811),
    .X(_06559_));
 sky130_fd_sc_hd__mux4_1 _12848_ (.A0(\dpath.RF.R[0][21] ),
    .A1(\dpath.RF.R[1][21] ),
    .A2(\dpath.RF.R[2][21] ),
    .A3(\dpath.RF.R[3][21] ),
    .S0(net835),
    .S1(net811),
    .X(_06560_));
 sky130_fd_sc_hd__mux4_1 _12849_ (.A0(\dpath.RF.R[4][21] ),
    .A1(\dpath.RF.R[5][21] ),
    .A2(\dpath.RF.R[6][21] ),
    .A3(\dpath.RF.R[7][21] ),
    .S0(net835),
    .S1(net811),
    .X(_06561_));
 sky130_fd_sc_hd__mux4_1 _12850_ (.A0(_06558_),
    .A1(_06559_),
    .A2(_06561_),
    .A3(_06560_),
    .S0(net499),
    .S1(net493),
    .X(_06562_));
 sky130_fd_sc_hd__or2_1 _12851_ (.A(net792),
    .B(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__and3_1 _12852_ (.A(net363),
    .B(_06557_),
    .C(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__a22o_1 _12853_ (.A1(net676),
    .A2(net379),
    .B1(net357),
    .B2(_04003_),
    .X(_06565_));
 sky130_fd_sc_hd__a21o_1 _12854_ (.A1(_04113_),
    .A2(net377),
    .B1(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__a21oi_4 _12855_ (.A1(net359),
    .A2(_06566_),
    .B1(_06564_),
    .Y(_06567_));
 sky130_fd_sc_hd__o21a_1 _12856_ (.A1(net477),
    .A2(_06567_),
    .B1(net472),
    .X(_06568_));
 sky130_fd_sc_hd__nor2_1 _12857_ (.A(net885),
    .B(_06568_),
    .Y(_01174_));
 sky130_fd_sc_hd__mux4_1 _12858_ (.A0(\dpath.RF.R[24][22] ),
    .A1(\dpath.RF.R[25][22] ),
    .A2(\dpath.RF.R[26][22] ),
    .A3(\dpath.RF.R[27][22] ),
    .S0(net837),
    .S1(net814),
    .X(_06569_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(\dpath.RF.R[30][22] ),
    .A1(\dpath.RF.R[31][22] ),
    .S(net837),
    .X(_06570_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(\dpath.RF.R[28][22] ),
    .A1(\dpath.RF.R[29][22] ),
    .S(net837),
    .X(_06571_));
 sky130_fd_sc_hd__a21o_1 _12861_ (.A1(net504),
    .A2(_06571_),
    .B1(net500),
    .X(_06572_));
 sky130_fd_sc_hd__a21o_1 _12862_ (.A1(net814),
    .A2(_06570_),
    .B1(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__o211a_1 _12863_ (.A1(net798),
    .A2(_06569_),
    .B1(_06573_),
    .C1(net795),
    .X(_06574_));
 sky130_fd_sc_hd__mux4_1 _12864_ (.A0(\dpath.RF.R[20][22] ),
    .A1(\dpath.RF.R[21][22] ),
    .A2(\dpath.RF.R[22][22] ),
    .A3(\dpath.RF.R[23][22] ),
    .S0(net836),
    .S1(net814),
    .X(_06575_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(\dpath.RF.R[18][22] ),
    .A1(\dpath.RF.R[19][22] ),
    .S(net836),
    .X(_06576_));
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(\dpath.RF.R[16][22] ),
    .A1(\dpath.RF.R[17][22] ),
    .S(net836),
    .X(_06577_));
 sky130_fd_sc_hd__a21o_1 _12867_ (.A1(_01788_),
    .A2(_06577_),
    .B1(_00002_),
    .X(_06578_));
 sky130_fd_sc_hd__a21o_1 _12868_ (.A1(net814),
    .A2(_06576_),
    .B1(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__o211a_1 _12869_ (.A1(net500),
    .A2(_06575_),
    .B1(_06579_),
    .C1(_01790_),
    .X(_06580_));
 sky130_fd_sc_hd__or3b_1 _12870_ (.A(_06574_),
    .B(_06580_),
    .C_N(net793),
    .X(_06581_));
 sky130_fd_sc_hd__mux4_1 _12871_ (.A0(\dpath.RF.R[12][22] ),
    .A1(\dpath.RF.R[13][22] ),
    .A2(\dpath.RF.R[14][22] ),
    .A3(\dpath.RF.R[15][22] ),
    .S0(net836),
    .S1(net814),
    .X(_06582_));
 sky130_fd_sc_hd__mux4_1 _12872_ (.A0(\dpath.RF.R[8][22] ),
    .A1(\dpath.RF.R[9][22] ),
    .A2(\dpath.RF.R[10][22] ),
    .A3(\dpath.RF.R[11][22] ),
    .S0(net831),
    .S1(net810),
    .X(_06583_));
 sky130_fd_sc_hd__mux4_1 _12873_ (.A0(\dpath.RF.R[0][22] ),
    .A1(\dpath.RF.R[1][22] ),
    .A2(\dpath.RF.R[2][22] ),
    .A3(\dpath.RF.R[3][22] ),
    .S0(net836),
    .S1(net814),
    .X(_06584_));
 sky130_fd_sc_hd__mux4_1 _12874_ (.A0(\dpath.RF.R[4][22] ),
    .A1(\dpath.RF.R[5][22] ),
    .A2(\dpath.RF.R[6][22] ),
    .A3(\dpath.RF.R[7][22] ),
    .S0(net836),
    .S1(net814),
    .X(_06585_));
 sky130_fd_sc_hd__mux4_1 _12875_ (.A0(_06582_),
    .A1(_06583_),
    .A2(_06585_),
    .A3(_06584_),
    .S0(net500),
    .S1(net494),
    .X(_06586_));
 sky130_fd_sc_hd__or2_1 _12876_ (.A(net793),
    .B(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__and3_1 _12877_ (.A(net363),
    .B(_06581_),
    .C(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__a22o_1 _12878_ (.A1(net673),
    .A2(net379),
    .B1(net357),
    .B2(_04151_),
    .X(_06589_));
 sky130_fd_sc_hd__a21o_1 _12879_ (.A1(_04275_),
    .A2(net377),
    .B1(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__a21oi_4 _12880_ (.A1(net359),
    .A2(_06590_),
    .B1(_06588_),
    .Y(_06591_));
 sky130_fd_sc_hd__o21a_1 _12881_ (.A1(net477),
    .A2(_06591_),
    .B1(net472),
    .X(_06592_));
 sky130_fd_sc_hd__nor2_1 _12882_ (.A(net886),
    .B(_06592_),
    .Y(_01175_));
 sky130_fd_sc_hd__mux4_1 _12883_ (.A0(\dpath.RF.R[24][23] ),
    .A1(\dpath.RF.R[25][23] ),
    .A2(\dpath.RF.R[26][23] ),
    .A3(\dpath.RF.R[27][23] ),
    .S0(net838),
    .S1(net816),
    .X(_06593_));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(\dpath.RF.R[30][23] ),
    .A1(\dpath.RF.R[31][23] ),
    .S(net838),
    .X(_06594_));
 sky130_fd_sc_hd__mux2_1 _12885_ (.A0(\dpath.RF.R[28][23] ),
    .A1(\dpath.RF.R[29][23] ),
    .S(net838),
    .X(_06595_));
 sky130_fd_sc_hd__a21o_1 _12886_ (.A1(net504),
    .A2(_06595_),
    .B1(net501),
    .X(_06596_));
 sky130_fd_sc_hd__a21o_1 _12887_ (.A1(net816),
    .A2(_06594_),
    .B1(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__o211a_1 _12888_ (.A1(net798),
    .A2(_06593_),
    .B1(_06597_),
    .C1(net795),
    .X(_06598_));
 sky130_fd_sc_hd__mux4_1 _12889_ (.A0(\dpath.RF.R[20][23] ),
    .A1(\dpath.RF.R[21][23] ),
    .A2(\dpath.RF.R[22][23] ),
    .A3(\dpath.RF.R[23][23] ),
    .S0(net837),
    .S1(net814),
    .X(_06599_));
 sky130_fd_sc_hd__mux2_1 _12890_ (.A0(\dpath.RF.R[18][23] ),
    .A1(\dpath.RF.R[19][23] ),
    .S(net838),
    .X(_06600_));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(\dpath.RF.R[16][23] ),
    .A1(\dpath.RF.R[17][23] ),
    .S(net838),
    .X(_06601_));
 sky130_fd_sc_hd__a21o_1 _12892_ (.A1(net505),
    .A2(_06601_),
    .B1(_00002_),
    .X(_06602_));
 sky130_fd_sc_hd__a21o_1 _12893_ (.A1(net816),
    .A2(_06600_),
    .B1(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__o211a_1 _12894_ (.A1(net501),
    .A2(_06599_),
    .B1(_06603_),
    .C1(net494),
    .X(_06604_));
 sky130_fd_sc_hd__or3b_1 _12895_ (.A(_06598_),
    .B(_06604_),
    .C_N(net3665),
    .X(_06605_));
 sky130_fd_sc_hd__mux4_1 _12896_ (.A0(\dpath.RF.R[12][23] ),
    .A1(\dpath.RF.R[13][23] ),
    .A2(\dpath.RF.R[14][23] ),
    .A3(\dpath.RF.R[15][23] ),
    .S0(net834),
    .S1(net812),
    .X(_06606_));
 sky130_fd_sc_hd__mux4_1 _12897_ (.A0(\dpath.RF.R[8][23] ),
    .A1(\dpath.RF.R[9][23] ),
    .A2(\dpath.RF.R[10][23] ),
    .A3(\dpath.RF.R[11][23] ),
    .S0(net834),
    .S1(net812),
    .X(_06607_));
 sky130_fd_sc_hd__mux4_1 _12898_ (.A0(\dpath.RF.R[0][23] ),
    .A1(\dpath.RF.R[1][23] ),
    .A2(\dpath.RF.R[2][23] ),
    .A3(\dpath.RF.R[3][23] ),
    .S0(net831),
    .S1(net810),
    .X(_06608_));
 sky130_fd_sc_hd__mux4_1 _12899_ (.A0(\dpath.RF.R[4][23] ),
    .A1(\dpath.RF.R[5][23] ),
    .A2(\dpath.RF.R[6][23] ),
    .A3(\dpath.RF.R[7][23] ),
    .S0(net831),
    .S1(net810),
    .X(_06609_));
 sky130_fd_sc_hd__mux4_1 _12900_ (.A0(_06606_),
    .A1(_06607_),
    .A2(_06609_),
    .A3(_06608_),
    .S0(net499),
    .S1(net493),
    .X(_06610_));
 sky130_fd_sc_hd__or2_1 _12901_ (.A(net792),
    .B(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__and3_1 _12902_ (.A(net363),
    .B(_06605_),
    .C(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__a22o_1 _12903_ (.A1(net671),
    .A2(net379),
    .B1(net357),
    .B2(_04301_),
    .X(_06613_));
 sky130_fd_sc_hd__a21o_1 _12904_ (.A1(_04421_),
    .A2(net377),
    .B1(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__a21oi_4 _12905_ (.A1(net359),
    .A2(_06614_),
    .B1(_06612_),
    .Y(_06615_));
 sky130_fd_sc_hd__o21a_1 _12906_ (.A1(net477),
    .A2(_06615_),
    .B1(net472),
    .X(_06616_));
 sky130_fd_sc_hd__nor2_1 _12907_ (.A(net885),
    .B(_06616_),
    .Y(_01176_));
 sky130_fd_sc_hd__mux4_1 _12908_ (.A0(net3695),
    .A1(\dpath.RF.R[25][24] ),
    .A2(\dpath.RF.R[26][24] ),
    .A3(\dpath.RF.R[27][24] ),
    .S0(net834),
    .S1(net812),
    .X(_06617_));
 sky130_fd_sc_hd__mux2_1 _12909_ (.A0(net1250),
    .A1(\dpath.RF.R[31][24] ),
    .S(net835),
    .X(_06618_));
 sky130_fd_sc_hd__mux2_1 _12910_ (.A0(\dpath.RF.R[28][24] ),
    .A1(\dpath.RF.R[29][24] ),
    .S(net835),
    .X(_06619_));
 sky130_fd_sc_hd__a21o_1 _12911_ (.A1(net504),
    .A2(_06619_),
    .B1(net499),
    .X(_06620_));
 sky130_fd_sc_hd__a21o_1 _12912_ (.A1(net812),
    .A2(_06618_),
    .B1(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__o211a_1 _12913_ (.A1(net798),
    .A2(_06617_),
    .B1(_06621_),
    .C1(net795),
    .X(_06622_));
 sky130_fd_sc_hd__mux4_1 _12914_ (.A0(\dpath.RF.R[20][24] ),
    .A1(\dpath.RF.R[21][24] ),
    .A2(\dpath.RF.R[22][24] ),
    .A3(\dpath.RF.R[23][24] ),
    .S0(net834),
    .S1(net812),
    .X(_06623_));
 sky130_fd_sc_hd__mux2_1 _12915_ (.A0(\dpath.RF.R[18][24] ),
    .A1(\dpath.RF.R[19][24] ),
    .S(net835),
    .X(_06624_));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(\dpath.RF.R[16][24] ),
    .A1(\dpath.RF.R[17][24] ),
    .S(net834),
    .X(_06625_));
 sky130_fd_sc_hd__a21o_1 _12917_ (.A1(net504),
    .A2(_06625_),
    .B1(net798),
    .X(_06626_));
 sky130_fd_sc_hd__a21o_1 _12918_ (.A1(net813),
    .A2(_06624_),
    .B1(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__o211a_1 _12919_ (.A1(net499),
    .A2(_06623_),
    .B1(_06627_),
    .C1(net493),
    .X(_06628_));
 sky130_fd_sc_hd__or3b_1 _12920_ (.A(_06622_),
    .B(_06628_),
    .C_N(net792),
    .X(_06629_));
 sky130_fd_sc_hd__mux4_1 _12921_ (.A0(\dpath.RF.R[12][24] ),
    .A1(\dpath.RF.R[13][24] ),
    .A2(\dpath.RF.R[14][24] ),
    .A3(\dpath.RF.R[15][24] ),
    .S0(net834),
    .S1(net812),
    .X(_06630_));
 sky130_fd_sc_hd__mux4_1 _12922_ (.A0(\dpath.RF.R[8][24] ),
    .A1(\dpath.RF.R[9][24] ),
    .A2(\dpath.RF.R[10][24] ),
    .A3(\dpath.RF.R[11][24] ),
    .S0(net834),
    .S1(net812),
    .X(_06631_));
 sky130_fd_sc_hd__mux4_1 _12923_ (.A0(net1174),
    .A1(\dpath.RF.R[1][24] ),
    .A2(\dpath.RF.R[2][24] ),
    .A3(\dpath.RF.R[3][24] ),
    .S0(net834),
    .S1(net812),
    .X(_06632_));
 sky130_fd_sc_hd__mux4_1 _12924_ (.A0(\dpath.RF.R[4][24] ),
    .A1(\dpath.RF.R[5][24] ),
    .A2(\dpath.RF.R[6][24] ),
    .A3(\dpath.RF.R[7][24] ),
    .S0(net834),
    .S1(net812),
    .X(_06633_));
 sky130_fd_sc_hd__mux4_1 _12925_ (.A0(_06630_),
    .A1(_06631_),
    .A2(_06633_),
    .A3(_06632_),
    .S0(net499),
    .S1(net493),
    .X(_06634_));
 sky130_fd_sc_hd__or2_1 _12926_ (.A(net793),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__and3_1 _12927_ (.A(net363),
    .B(_06629_),
    .C(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__a22o_1 _12928_ (.A1(net670),
    .A2(net379),
    .B1(net357),
    .B2(_04452_),
    .X(_06637_));
 sky130_fd_sc_hd__a21o_1 _12929_ (.A1(_04593_),
    .A2(net377),
    .B1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__a21oi_4 _12930_ (.A1(net359),
    .A2(_06638_),
    .B1(_06636_),
    .Y(_06639_));
 sky130_fd_sc_hd__o21a_1 _12931_ (.A1(net477),
    .A2(_06639_),
    .B1(net472),
    .X(_06640_));
 sky130_fd_sc_hd__nor2_1 _12932_ (.A(net885),
    .B(_06640_),
    .Y(_01177_));
 sky130_fd_sc_hd__mux4_1 _12933_ (.A0(\dpath.RF.R[24][25] ),
    .A1(\dpath.RF.R[25][25] ),
    .A2(\dpath.RF.R[26][25] ),
    .A3(\dpath.RF.R[27][25] ),
    .S0(net834),
    .S1(net812),
    .X(_06641_));
 sky130_fd_sc_hd__mux2_1 _12934_ (.A0(\dpath.RF.R[30][25] ),
    .A1(\dpath.RF.R[31][25] ),
    .S(net838),
    .X(_06642_));
 sky130_fd_sc_hd__mux2_1 _12935_ (.A0(\dpath.RF.R[28][25] ),
    .A1(\dpath.RF.R[29][25] ),
    .S(net838),
    .X(_06643_));
 sky130_fd_sc_hd__a21o_1 _12936_ (.A1(net505),
    .A2(_06643_),
    .B1(net501),
    .X(_06644_));
 sky130_fd_sc_hd__a21o_1 _12937_ (.A1(net816),
    .A2(_06642_),
    .B1(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__o211a_1 _12938_ (.A1(net799),
    .A2(_06641_),
    .B1(_06645_),
    .C1(net795),
    .X(_06646_));
 sky130_fd_sc_hd__mux4_1 _12939_ (.A0(\dpath.RF.R[20][25] ),
    .A1(\dpath.RF.R[21][25] ),
    .A2(\dpath.RF.R[22][25] ),
    .A3(\dpath.RF.R[23][25] ),
    .S0(net835),
    .S1(net813),
    .X(_06647_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(\dpath.RF.R[18][25] ),
    .A1(\dpath.RF.R[19][25] ),
    .S(net838),
    .X(_06648_));
 sky130_fd_sc_hd__mux2_1 _12941_ (.A0(\dpath.RF.R[16][25] ),
    .A1(\dpath.RF.R[17][25] ),
    .S(net838),
    .X(_06649_));
 sky130_fd_sc_hd__a21o_1 _12942_ (.A1(net505),
    .A2(_06649_),
    .B1(net799),
    .X(_06650_));
 sky130_fd_sc_hd__a21o_1 _12943_ (.A1(net818),
    .A2(_06648_),
    .B1(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__o211a_1 _12944_ (.A1(net499),
    .A2(_06647_),
    .B1(_06651_),
    .C1(net493),
    .X(_06652_));
 sky130_fd_sc_hd__or3b_1 _12945_ (.A(_06646_),
    .B(_06652_),
    .C_N(net793),
    .X(_06653_));
 sky130_fd_sc_hd__mux4_1 _12946_ (.A0(\dpath.RF.R[12][25] ),
    .A1(\dpath.RF.R[13][25] ),
    .A2(\dpath.RF.R[14][25] ),
    .A3(\dpath.RF.R[15][25] ),
    .S0(net838),
    .S1(net816),
    .X(_06654_));
 sky130_fd_sc_hd__mux4_1 _12947_ (.A0(\dpath.RF.R[8][25] ),
    .A1(\dpath.RF.R[9][25] ),
    .A2(\dpath.RF.R[10][25] ),
    .A3(\dpath.RF.R[11][25] ),
    .S0(net839),
    .S1(net818),
    .X(_06655_));
 sky130_fd_sc_hd__mux4_1 _12948_ (.A0(\dpath.RF.R[0][25] ),
    .A1(\dpath.RF.R[1][25] ),
    .A2(\dpath.RF.R[2][25] ),
    .A3(\dpath.RF.R[3][25] ),
    .S0(net834),
    .S1(net812),
    .X(_06656_));
 sky130_fd_sc_hd__mux4_1 _12949_ (.A0(\dpath.RF.R[4][25] ),
    .A1(\dpath.RF.R[5][25] ),
    .A2(\dpath.RF.R[6][25] ),
    .A3(\dpath.RF.R[7][25] ),
    .S0(net835),
    .S1(net812),
    .X(_06657_));
 sky130_fd_sc_hd__mux4_1 _12950_ (.A0(_06654_),
    .A1(_06655_),
    .A2(_06657_),
    .A3(_06656_),
    .S0(net499),
    .S1(net494),
    .X(_06658_));
 sky130_fd_sc_hd__or2_1 _12951_ (.A(net792),
    .B(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__and3_1 _12952_ (.A(net363),
    .B(_06653_),
    .C(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__a22o_1 _12953_ (.A1(net667),
    .A2(net380),
    .B1(net358),
    .B2(_04627_),
    .X(_06661_));
 sky130_fd_sc_hd__a21o_1 _12954_ (.A1(_04759_),
    .A2(net378),
    .B1(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__a21oi_2 _12955_ (.A1(net360),
    .A2(_06662_),
    .B1(_06660_),
    .Y(_06663_));
 sky130_fd_sc_hd__o21a_1 _12956_ (.A1(net477),
    .A2(_06663_),
    .B1(net472),
    .X(_06664_));
 sky130_fd_sc_hd__nor2_1 _12957_ (.A(net885),
    .B(_06664_),
    .Y(_01178_));
 sky130_fd_sc_hd__mux4_1 _12958_ (.A0(net1714),
    .A1(net1722),
    .A2(net2428),
    .A3(net2930),
    .S0(net842),
    .S1(net815),
    .X(_06665_));
 sky130_fd_sc_hd__mux2_1 _12959_ (.A0(net1728),
    .A1(net3106),
    .S(net837),
    .X(_06666_));
 sky130_fd_sc_hd__mux2_1 _12960_ (.A0(net2568),
    .A1(net2466),
    .S(net837),
    .X(_06667_));
 sky130_fd_sc_hd__a21o_1 _12961_ (.A1(net505),
    .A2(_06667_),
    .B1(net500),
    .X(_06668_));
 sky130_fd_sc_hd__a21o_1 _12962_ (.A1(net815),
    .A2(_06666_),
    .B1(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__o211a_1 _12963_ (.A1(net799),
    .A2(_06665_),
    .B1(_06669_),
    .C1(net795),
    .X(_06670_));
 sky130_fd_sc_hd__mux4_1 _12964_ (.A0(net2732),
    .A1(net2516),
    .A2(net2494),
    .A3(net3196),
    .S0(net842),
    .S1(net815),
    .X(_06671_));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(net3108),
    .A1(net1902),
    .S(net837),
    .X(_06672_));
 sky130_fd_sc_hd__mux2_1 _12966_ (.A0(\dpath.RF.R[16][26] ),
    .A1(net1328),
    .S(net837),
    .X(_06673_));
 sky130_fd_sc_hd__a21o_1 _12967_ (.A1(net505),
    .A2(_06673_),
    .B1(net799),
    .X(_06674_));
 sky130_fd_sc_hd__a21o_1 _12968_ (.A1(net815),
    .A2(_06672_),
    .B1(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__o211a_1 _12969_ (.A1(net500),
    .A2(_06671_),
    .B1(_06675_),
    .C1(net494),
    .X(_06676_));
 sky130_fd_sc_hd__or3b_1 _12970_ (.A(_06670_),
    .B(_06676_),
    .C_N(net793),
    .X(_06677_));
 sky130_fd_sc_hd__mux4_1 _12971_ (.A0(\dpath.RF.R[12][26] ),
    .A1(net1344),
    .A2(\dpath.RF.R[14][26] ),
    .A3(net2676),
    .S0(net836),
    .S1(net814),
    .X(_06678_));
 sky130_fd_sc_hd__mux4_1 _12972_ (.A0(\dpath.RF.R[8][26] ),
    .A1(\dpath.RF.R[9][26] ),
    .A2(\dpath.RF.R[10][26] ),
    .A3(\dpath.RF.R[11][26] ),
    .S0(net836),
    .S1(net814),
    .X(_06679_));
 sky130_fd_sc_hd__mux4_1 _12973_ (.A0(\dpath.RF.R[0][26] ),
    .A1(\dpath.RF.R[1][26] ),
    .A2(net2140),
    .A3(\dpath.RF.R[3][26] ),
    .S0(net836),
    .S1(net814),
    .X(_06680_));
 sky130_fd_sc_hd__mux4_1 _12974_ (.A0(\dpath.RF.R[4][26] ),
    .A1(\dpath.RF.R[5][26] ),
    .A2(\dpath.RF.R[6][26] ),
    .A3(\dpath.RF.R[7][26] ),
    .S0(net836),
    .S1(net814),
    .X(_06681_));
 sky130_fd_sc_hd__mux4_1 _12975_ (.A0(_06678_),
    .A1(_06679_),
    .A2(_06681_),
    .A3(_06680_),
    .S0(net500),
    .S1(net494),
    .X(_06682_));
 sky130_fd_sc_hd__or2_1 _12976_ (.A(net793),
    .B(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__and3_1 _12977_ (.A(net363),
    .B(_06677_),
    .C(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__a22o_1 _12978_ (.A1(net3660),
    .A2(net379),
    .B1(net357),
    .B2(_04789_),
    .X(_06685_));
 sky130_fd_sc_hd__a21o_1 _12979_ (.A1(_04933_),
    .A2(net377),
    .B1(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__a21oi_1 _12980_ (.A1(net359),
    .A2(_06686_),
    .B1(_06684_),
    .Y(_06687_));
 sky130_fd_sc_hd__o21a_1 _12981_ (.A1(net477),
    .A2(_06687_),
    .B1(_02844_),
    .X(_06688_));
 sky130_fd_sc_hd__nor2_1 _12982_ (.A(net886),
    .B(_06688_),
    .Y(_01179_));
 sky130_fd_sc_hd__mux4_1 _12983_ (.A0(net2554),
    .A1(net1764),
    .A2(net1932),
    .A3(net1668),
    .S0(net838),
    .S1(net816),
    .X(_06689_));
 sky130_fd_sc_hd__mux2_1 _12984_ (.A0(net1610),
    .A1(net3144),
    .S(net839),
    .X(_06690_));
 sky130_fd_sc_hd__mux2_1 _12985_ (.A0(net2668),
    .A1(net3128),
    .S(net839),
    .X(_06691_));
 sky130_fd_sc_hd__a21o_1 _12986_ (.A1(net505),
    .A2(_06691_),
    .B1(net501),
    .X(_06692_));
 sky130_fd_sc_hd__a21o_1 _12987_ (.A1(net816),
    .A2(_06690_),
    .B1(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__o211a_1 _12988_ (.A1(net799),
    .A2(_06689_),
    .B1(_06693_),
    .C1(net795),
    .X(_06694_));
 sky130_fd_sc_hd__mux4_1 _12989_ (.A0(net2756),
    .A1(net2492),
    .A2(net1528),
    .A3(net2408),
    .S0(net838),
    .S1(net816),
    .X(_06695_));
 sky130_fd_sc_hd__mux2_1 _12990_ (.A0(net1204),
    .A1(net1654),
    .S(net839),
    .X(_06696_));
 sky130_fd_sc_hd__mux2_1 _12991_ (.A0(net1630),
    .A1(net1798),
    .S(net839),
    .X(_06697_));
 sky130_fd_sc_hd__a21o_1 _12992_ (.A1(net505),
    .A2(_06697_),
    .B1(net799),
    .X(_06698_));
 sky130_fd_sc_hd__a21o_1 _12993_ (.A1(net816),
    .A2(_06696_),
    .B1(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__o211a_1 _12994_ (.A1(net501),
    .A2(_06695_),
    .B1(_06699_),
    .C1(net494),
    .X(_06700_));
 sky130_fd_sc_hd__or3b_1 _12995_ (.A(_06694_),
    .B(_06700_),
    .C_N(net793),
    .X(_06701_));
 sky130_fd_sc_hd__mux4_1 _12996_ (.A0(net2260),
    .A1(net2504),
    .A2(net1448),
    .A3(net2862),
    .S0(net838),
    .S1(net816),
    .X(_06702_));
 sky130_fd_sc_hd__mux4_1 _12997_ (.A0(net1458),
    .A1(net1744),
    .A2(net1376),
    .A3(net2000),
    .S0(net839),
    .S1(net816),
    .X(_06703_));
 sky130_fd_sc_hd__mux4_1 _12998_ (.A0(net1052),
    .A1(net2778),
    .A2(net1518),
    .A3(net2072),
    .S0(net839),
    .S1(net816),
    .X(_06704_));
 sky130_fd_sc_hd__mux4_1 _12999_ (.A0(net2232),
    .A1(net1670),
    .A2(net2582),
    .A3(net3130),
    .S0(net839),
    .S1(net816),
    .X(_06705_));
 sky130_fd_sc_hd__mux4_1 _13000_ (.A0(_06702_),
    .A1(_06703_),
    .A2(_06705_),
    .A3(_06704_),
    .S0(net501),
    .S1(net494),
    .X(_06706_));
 sky130_fd_sc_hd__or2_1 _13001_ (.A(net793),
    .B(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__and3_1 _13002_ (.A(net363),
    .B(_06701_),
    .C(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__a22o_1 _13003_ (.A1(net663),
    .A2(net379),
    .B1(net357),
    .B2(_04968_),
    .X(_06709_));
 sky130_fd_sc_hd__a21o_1 _13004_ (.A1(_05109_),
    .A2(net377),
    .B1(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a21oi_2 _13005_ (.A1(net359),
    .A2(_06710_),
    .B1(_06708_),
    .Y(_06711_));
 sky130_fd_sc_hd__o21a_1 _13006_ (.A1(net478),
    .A2(_06711_),
    .B1(net472),
    .X(_06712_));
 sky130_fd_sc_hd__nor2_1 _13007_ (.A(net885),
    .B(_06712_),
    .Y(_01180_));
 sky130_fd_sc_hd__mux4_1 _13008_ (.A0(net1702),
    .A1(net2386),
    .A2(net1626),
    .A3(net2524),
    .S0(net840),
    .S1(net817),
    .X(_06713_));
 sky130_fd_sc_hd__mux2_1 _13009_ (.A0(net1470),
    .A1(net3030),
    .S(net840),
    .X(_06714_));
 sky130_fd_sc_hd__mux2_1 _13010_ (.A0(net1546),
    .A1(net2852),
    .S(net840),
    .X(_06715_));
 sky130_fd_sc_hd__a21o_1 _13011_ (.A1(net505),
    .A2(_06715_),
    .B1(net500),
    .X(_06716_));
 sky130_fd_sc_hd__a21o_1 _13012_ (.A1(net817),
    .A2(_06714_),
    .B1(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__o211a_1 _13013_ (.A1(net799),
    .A2(_06713_),
    .B1(_06717_),
    .C1(net3669),
    .X(_06718_));
 sky130_fd_sc_hd__mux4_1 _13014_ (.A0(net1494),
    .A1(net1730),
    .A2(net1388),
    .A3(net1894),
    .S0(net840),
    .S1(net817),
    .X(_06719_));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(net1974),
    .A1(net2520),
    .S(net840),
    .X(_06720_));
 sky130_fd_sc_hd__mux2_1 _13016_ (.A0(net1990),
    .A1(net1562),
    .S(net840),
    .X(_06721_));
 sky130_fd_sc_hd__a21o_1 _13017_ (.A1(net505),
    .A2(_06721_),
    .B1(net799),
    .X(_06722_));
 sky130_fd_sc_hd__a21o_1 _13018_ (.A1(net817),
    .A2(_06720_),
    .B1(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__o211a_1 _13019_ (.A1(net500),
    .A2(_06719_),
    .B1(_06723_),
    .C1(net494),
    .X(_06724_));
 sky130_fd_sc_hd__or3b_1 _13020_ (.A(_06718_),
    .B(_06724_),
    .C_N(net793),
    .X(_06725_));
 sky130_fd_sc_hd__mux4_1 _13021_ (.A0(net2496),
    .A1(net1858),
    .A2(net1306),
    .A3(net2430),
    .S0(net840),
    .S1(net817),
    .X(_06726_));
 sky130_fd_sc_hd__mux4_1 _13022_ (.A0(net1266),
    .A1(net1244),
    .A2(net1258),
    .A3(net2904),
    .S0(net838),
    .S1(net816),
    .X(_06727_));
 sky130_fd_sc_hd__mux4_1 _13023_ (.A0(net1154),
    .A1(\dpath.RF.R[1][28] ),
    .A2(net1598),
    .A3(\dpath.RF.R[3][28] ),
    .S0(net838),
    .S1(net816),
    .X(_06728_));
 sky130_fd_sc_hd__mux4_1 _13024_ (.A0(\dpath.RF.R[4][28] ),
    .A1(\dpath.RF.R[5][28] ),
    .A2(\dpath.RF.R[6][28] ),
    .A3(\dpath.RF.R[7][28] ),
    .S0(net838),
    .S1(net816),
    .X(_06729_));
 sky130_fd_sc_hd__mux4_1 _13025_ (.A0(_06726_),
    .A1(_06727_),
    .A2(_06729_),
    .A3(_06728_),
    .S0(net501),
    .S1(net494),
    .X(_06730_));
 sky130_fd_sc_hd__or2_1 _13026_ (.A(net793),
    .B(_06730_),
    .X(_06731_));
 sky130_fd_sc_hd__and3_1 _13027_ (.A(net364),
    .B(net3670),
    .C(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__a22o_1 _13028_ (.A1(net661),
    .A2(net380),
    .B1(net357),
    .B2(_05139_),
    .X(_06733_));
 sky130_fd_sc_hd__a21o_1 _13029_ (.A1(_05292_),
    .A2(net377),
    .B1(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__a21oi_2 _13030_ (.A1(net359),
    .A2(_06734_),
    .B1(net3671),
    .Y(_06735_));
 sky130_fd_sc_hd__o21a_1 _13031_ (.A1(_01975_),
    .A2(_06735_),
    .B1(net472),
    .X(_06736_));
 sky130_fd_sc_hd__nor2_1 _13032_ (.A(net886),
    .B(_06736_),
    .Y(_01181_));
 sky130_fd_sc_hd__mux4_1 _13033_ (.A0(\dpath.RF.R[24][29] ),
    .A1(\dpath.RF.R[25][29] ),
    .A2(\dpath.RF.R[26][29] ),
    .A3(\dpath.RF.R[27][29] ),
    .S0(net840),
    .S1(net817),
    .X(_06737_));
 sky130_fd_sc_hd__mux2_1 _13034_ (.A0(\dpath.RF.R[30][29] ),
    .A1(\dpath.RF.R[31][29] ),
    .S(net840),
    .X(_06738_));
 sky130_fd_sc_hd__mux2_1 _13035_ (.A0(\dpath.RF.R[28][29] ),
    .A1(\dpath.RF.R[29][29] ),
    .S(net840),
    .X(_06739_));
 sky130_fd_sc_hd__a21o_1 _13036_ (.A1(net505),
    .A2(_06739_),
    .B1(net500),
    .X(_06740_));
 sky130_fd_sc_hd__a21o_1 _13037_ (.A1(net817),
    .A2(_06738_),
    .B1(_06740_),
    .X(_06741_));
 sky130_fd_sc_hd__o211a_1 _13038_ (.A1(net799),
    .A2(_06737_),
    .B1(_06741_),
    .C1(net3669),
    .X(_06742_));
 sky130_fd_sc_hd__mux4_1 _13039_ (.A0(net1708),
    .A1(\dpath.RF.R[21][29] ),
    .A2(\dpath.RF.R[22][29] ),
    .A3(\dpath.RF.R[23][29] ),
    .S0(net840),
    .S1(net817),
    .X(_06743_));
 sky130_fd_sc_hd__mux2_1 _13040_ (.A0(net1384),
    .A1(net2134),
    .S(net841),
    .X(_06744_));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(\dpath.RF.R[16][29] ),
    .A1(\dpath.RF.R[17][29] ),
    .S(net840),
    .X(_06745_));
 sky130_fd_sc_hd__a21o_1 _13042_ (.A1(net505),
    .A2(_06745_),
    .B1(net799),
    .X(_06746_));
 sky130_fd_sc_hd__a21o_1 _13043_ (.A1(net818),
    .A2(_06744_),
    .B1(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__o211a_1 _13044_ (.A1(net500),
    .A2(_06743_),
    .B1(_06747_),
    .C1(net494),
    .X(_06748_));
 sky130_fd_sc_hd__or3b_1 _13045_ (.A(_06742_),
    .B(_06748_),
    .C_N(net793),
    .X(_06749_));
 sky130_fd_sc_hd__mux4_1 _13046_ (.A0(\dpath.RF.R[12][29] ),
    .A1(\dpath.RF.R[13][29] ),
    .A2(\dpath.RF.R[14][29] ),
    .A3(\dpath.RF.R[15][29] ),
    .S0(net841),
    .S1(net818),
    .X(_06750_));
 sky130_fd_sc_hd__mux4_1 _13047_ (.A0(\dpath.RF.R[8][29] ),
    .A1(\dpath.RF.R[9][29] ),
    .A2(\dpath.RF.R[10][29] ),
    .A3(\dpath.RF.R[11][29] ),
    .S0(net840),
    .S1(net817),
    .X(_06751_));
 sky130_fd_sc_hd__mux4_1 _13048_ (.A0(\dpath.RF.R[0][29] ),
    .A1(\dpath.RF.R[1][29] ),
    .A2(\dpath.RF.R[2][29] ),
    .A3(\dpath.RF.R[3][29] ),
    .S0(net841),
    .S1(net818),
    .X(_06752_));
 sky130_fd_sc_hd__mux4_1 _13049_ (.A0(\dpath.RF.R[4][29] ),
    .A1(\dpath.RF.R[5][29] ),
    .A2(\dpath.RF.R[6][29] ),
    .A3(\dpath.RF.R[7][29] ),
    .S0(net840),
    .S1(net817),
    .X(_06753_));
 sky130_fd_sc_hd__mux4_1 _13050_ (.A0(_06750_),
    .A1(_06751_),
    .A2(_06753_),
    .A3(_06752_),
    .S0(net501),
    .S1(net494),
    .X(_06754_));
 sky130_fd_sc_hd__or2_1 _13051_ (.A(net793),
    .B(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__and3_1 _13052_ (.A(net363),
    .B(_06749_),
    .C(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__a22o_1 _13053_ (.A1(net659),
    .A2(net379),
    .B1(net357),
    .B2(_05328_),
    .X(_06757_));
 sky130_fd_sc_hd__a21o_1 _13054_ (.A1(_05476_),
    .A2(net377),
    .B1(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__a21oi_1 _13055_ (.A1(net359),
    .A2(_06758_),
    .B1(_06756_),
    .Y(_06759_));
 sky130_fd_sc_hd__o21a_1 _13056_ (.A1(_01975_),
    .A2(_06759_),
    .B1(_02844_),
    .X(_06760_));
 sky130_fd_sc_hd__nor2_1 _13057_ (.A(net886),
    .B(_06760_),
    .Y(_01182_));
 sky130_fd_sc_hd__mux4_1 _13058_ (.A0(net1678),
    .A1(net2790),
    .A2(net1550),
    .A3(net1690),
    .S0(net837),
    .S1(net815),
    .X(_06761_));
 sky130_fd_sc_hd__mux2_1 _13059_ (.A0(net1294),
    .A1(\dpath.RF.R[31][30] ),
    .S(net837),
    .X(_06762_));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(\dpath.RF.R[28][30] ),
    .A1(\dpath.RF.R[29][30] ),
    .S(net837),
    .X(_06763_));
 sky130_fd_sc_hd__a21o_1 _13061_ (.A1(net505),
    .A2(_06763_),
    .B1(net500),
    .X(_06764_));
 sky130_fd_sc_hd__a21o_1 _13062_ (.A1(net815),
    .A2(_06762_),
    .B1(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__o211a_1 _13063_ (.A1(net799),
    .A2(_06761_),
    .B1(_06765_),
    .C1(_00003_),
    .X(_06766_));
 sky130_fd_sc_hd__mux4_1 _13064_ (.A0(net2324),
    .A1(net1718),
    .A2(net1252),
    .A3(net2288),
    .S0(net837),
    .S1(net815),
    .X(_06767_));
 sky130_fd_sc_hd__mux2_1 _13065_ (.A0(net1368),
    .A1(net2802),
    .S(net837),
    .X(_06768_));
 sky130_fd_sc_hd__mux2_1 _13066_ (.A0(\dpath.RF.R[16][30] ),
    .A1(\dpath.RF.R[17][30] ),
    .S(net837),
    .X(_06769_));
 sky130_fd_sc_hd__a21o_1 _13067_ (.A1(net505),
    .A2(_06769_),
    .B1(net799),
    .X(_06770_));
 sky130_fd_sc_hd__a21o_1 _13068_ (.A1(net815),
    .A2(_06768_),
    .B1(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__o211a_1 _13069_ (.A1(net500),
    .A2(_06767_),
    .B1(_06771_),
    .C1(net494),
    .X(_06772_));
 sky130_fd_sc_hd__or3b_1 _13070_ (.A(_06766_),
    .B(_06772_),
    .C_N(net793),
    .X(_06773_));
 sky130_fd_sc_hd__mux4_1 _13071_ (.A0(\dpath.RF.R[12][30] ),
    .A1(\dpath.RF.R[13][30] ),
    .A2(\dpath.RF.R[14][30] ),
    .A3(\dpath.RF.R[15][30] ),
    .S0(net836),
    .S1(net814),
    .X(_06774_));
 sky130_fd_sc_hd__mux4_1 _13072_ (.A0(\dpath.RF.R[8][30] ),
    .A1(\dpath.RF.R[9][30] ),
    .A2(\dpath.RF.R[10][30] ),
    .A3(\dpath.RF.R[11][30] ),
    .S0(net837),
    .S1(net814),
    .X(_06775_));
 sky130_fd_sc_hd__mux4_1 _13073_ (.A0(\dpath.RF.R[0][30] ),
    .A1(\dpath.RF.R[1][30] ),
    .A2(\dpath.RF.R[2][30] ),
    .A3(\dpath.RF.R[3][30] ),
    .S0(net836),
    .S1(net814),
    .X(_06776_));
 sky130_fd_sc_hd__mux4_1 _13074_ (.A0(\dpath.RF.R[4][30] ),
    .A1(\dpath.RF.R[5][30] ),
    .A2(\dpath.RF.R[6][30] ),
    .A3(\dpath.RF.R[7][30] ),
    .S0(net836),
    .S1(net814),
    .X(_06777_));
 sky130_fd_sc_hd__mux4_1 _13075_ (.A0(_06774_),
    .A1(_06775_),
    .A2(_06777_),
    .A3(_06776_),
    .S0(net500),
    .S1(net494),
    .X(_06778_));
 sky130_fd_sc_hd__or2_1 _13076_ (.A(net3665),
    .B(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__and3_1 _13077_ (.A(net363),
    .B(_06773_),
    .C(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__a22o_1 _13078_ (.A1(net656),
    .A2(net379),
    .B1(net357),
    .B2(_05509_),
    .X(_06781_));
 sky130_fd_sc_hd__a21o_1 _13079_ (.A1(_05662_),
    .A2(net377),
    .B1(_06781_),
    .X(_06782_));
 sky130_fd_sc_hd__a21oi_1 _13080_ (.A1(net359),
    .A2(_06782_),
    .B1(net3666),
    .Y(_06783_));
 sky130_fd_sc_hd__o21a_1 _13081_ (.A1(net478),
    .A2(_06783_),
    .B1(_02844_),
    .X(_06784_));
 sky130_fd_sc_hd__nor2_1 _13082_ (.A(net886),
    .B(_06784_),
    .Y(_01183_));
 sky130_fd_sc_hd__mux4_1 _13083_ (.A0(net2150),
    .A1(net2536),
    .A2(net1466),
    .A3(net2284),
    .S0(net840),
    .S1(net817),
    .X(_06785_));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(net1256),
    .A1(net2898),
    .S(net841),
    .X(_06786_));
 sky130_fd_sc_hd__mux2_1 _13085_ (.A0(\dpath.RF.R[28][31] ),
    .A1(\dpath.RF.R[29][31] ),
    .S(net841),
    .X(_06787_));
 sky130_fd_sc_hd__a21o_1 _13086_ (.A1(net505),
    .A2(_06787_),
    .B1(net500),
    .X(_06788_));
 sky130_fd_sc_hd__a21o_1 _13087_ (.A1(net817),
    .A2(_06786_),
    .B1(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__o211a_1 _13088_ (.A1(net799),
    .A2(_06785_),
    .B1(_06789_),
    .C1(net3669),
    .X(_06790_));
 sky130_fd_sc_hd__mux4_1 _13089_ (.A0(\dpath.RF.R[20][31] ),
    .A1(\dpath.RF.R[21][31] ),
    .A2(\dpath.RF.R[22][31] ),
    .A3(\dpath.RF.R[23][31] ),
    .S0(net840),
    .S1(net817),
    .X(_06791_));
 sky130_fd_sc_hd__mux2_1 _13090_ (.A0(\dpath.RF.R[18][31] ),
    .A1(\dpath.RF.R[19][31] ),
    .S(net841),
    .X(_06792_));
 sky130_fd_sc_hd__mux2_1 _13091_ (.A0(\dpath.RF.R[16][31] ),
    .A1(\dpath.RF.R[17][31] ),
    .S(net841),
    .X(_06793_));
 sky130_fd_sc_hd__a21o_1 _13092_ (.A1(net505),
    .A2(_06793_),
    .B1(net799),
    .X(_06794_));
 sky130_fd_sc_hd__a21o_1 _13093_ (.A1(net818),
    .A2(_06792_),
    .B1(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__o211a_1 _13094_ (.A1(net500),
    .A2(_06791_),
    .B1(_06795_),
    .C1(net494),
    .X(_06796_));
 sky130_fd_sc_hd__or3b_1 _13095_ (.A(_06790_),
    .B(_06796_),
    .C_N(net3665),
    .X(_06797_));
 sky130_fd_sc_hd__mux4_1 _13096_ (.A0(\dpath.RF.R[12][31] ),
    .A1(\dpath.RF.R[13][31] ),
    .A2(\dpath.RF.R[14][31] ),
    .A3(\dpath.RF.R[15][31] ),
    .S0(net841),
    .S1(net817),
    .X(_06798_));
 sky130_fd_sc_hd__mux4_1 _13097_ (.A0(\dpath.RF.R[8][31] ),
    .A1(\dpath.RF.R[9][31] ),
    .A2(\dpath.RF.R[10][31] ),
    .A3(\dpath.RF.R[11][31] ),
    .S0(net841),
    .S1(net817),
    .X(_06799_));
 sky130_fd_sc_hd__mux4_1 _13098_ (.A0(\dpath.RF.R[0][31] ),
    .A1(\dpath.RF.R[1][31] ),
    .A2(\dpath.RF.R[2][31] ),
    .A3(\dpath.RF.R[3][31] ),
    .S0(net841),
    .S1(net818),
    .X(_06800_));
 sky130_fd_sc_hd__mux4_1 _13099_ (.A0(\dpath.RF.R[4][31] ),
    .A1(\dpath.RF.R[5][31] ),
    .A2(\dpath.RF.R[6][31] ),
    .A3(\dpath.RF.R[7][31] ),
    .S0(net841),
    .S1(net817),
    .X(_06801_));
 sky130_fd_sc_hd__mux4_1 _13100_ (.A0(_06798_),
    .A1(_06799_),
    .A2(_06801_),
    .A3(_06800_),
    .S0(net500),
    .S1(net494),
    .X(_06802_));
 sky130_fd_sc_hd__or2_1 _13101_ (.A(net793),
    .B(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__and3_1 _13102_ (.A(net363),
    .B(_06797_),
    .C(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__a22o_1 _13103_ (.A1(net655),
    .A2(net379),
    .B1(_06063_),
    .B2(_05700_),
    .X(_06805_));
 sky130_fd_sc_hd__a21o_1 _13104_ (.A1(_05828_),
    .A2(net377),
    .B1(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__a21oi_1 _13105_ (.A1(net360),
    .A2(_06806_),
    .B1(_06804_),
    .Y(_06807_));
 sky130_fd_sc_hd__o21a_1 _13106_ (.A1(net477),
    .A2(_06807_),
    .B1(_02844_),
    .X(_06808_));
 sky130_fd_sc_hd__nor2_1 _13107_ (.A(net886),
    .B(_06808_),
    .Y(_01184_));
 sky130_fd_sc_hd__and2_1 _13108_ (.A(net874),
    .B(net958),
    .X(_01185_));
 sky130_fd_sc_hd__and2_1 _13109_ (.A(net873),
    .B(net1054),
    .X(_01186_));
 sky130_fd_sc_hd__and2_1 _13110_ (.A(net869),
    .B(net964),
    .X(_01187_));
 sky130_fd_sc_hd__and2_1 _13111_ (.A(net866),
    .B(net956),
    .X(_01188_));
 sky130_fd_sc_hd__and2_1 _13112_ (.A(net866),
    .B(net1010),
    .X(_01189_));
 sky130_fd_sc_hd__and2_1 _13113_ (.A(net866),
    .B(net940),
    .X(_01190_));
 sky130_fd_sc_hd__and2_1 _13114_ (.A(net867),
    .B(net946),
    .X(_01191_));
 sky130_fd_sc_hd__and2_1 _13115_ (.A(net869),
    .B(net950),
    .X(_01192_));
 sky130_fd_sc_hd__and2_1 _13116_ (.A(net870),
    .B(net916),
    .X(_01193_));
 sky130_fd_sc_hd__and2_1 _13117_ (.A(net869),
    .B(net926),
    .X(_01194_));
 sky130_fd_sc_hd__and2_1 _13118_ (.A(net870),
    .B(net976),
    .X(_01195_));
 sky130_fd_sc_hd__and2_1 _13119_ (.A(net866),
    .B(net962),
    .X(_01196_));
 sky130_fd_sc_hd__and2_1 _13120_ (.A(net868),
    .B(net1042),
    .X(_01197_));
 sky130_fd_sc_hd__and2_1 _13121_ (.A(net868),
    .B(net896),
    .X(_01198_));
 sky130_fd_sc_hd__and2_1 _13122_ (.A(net867),
    .B(net966),
    .X(_01199_));
 sky130_fd_sc_hd__and2_1 _13123_ (.A(net870),
    .B(net968),
    .X(_01200_));
 sky130_fd_sc_hd__and2_1 _13124_ (.A(net866),
    .B(net920),
    .X(_01201_));
 sky130_fd_sc_hd__and2_1 _13125_ (.A(net870),
    .B(net970),
    .X(_01202_));
 sky130_fd_sc_hd__and2_1 _13126_ (.A(net866),
    .B(net978),
    .X(_01203_));
 sky130_fd_sc_hd__and2_1 _13127_ (.A(net869),
    .B(net934),
    .X(_01204_));
 sky130_fd_sc_hd__and2_1 _13128_ (.A(net867),
    .B(net1032),
    .X(_01205_));
 sky130_fd_sc_hd__and2_1 _13129_ (.A(net866),
    .B(net988),
    .X(_01206_));
 sky130_fd_sc_hd__and2_1 _13130_ (.A(net869),
    .B(net928),
    .X(_01207_));
 sky130_fd_sc_hd__and2_1 _13131_ (.A(net873),
    .B(net1012),
    .X(_01208_));
 sky130_fd_sc_hd__and2_1 _13132_ (.A(net873),
    .B(net1048),
    .X(_01209_));
 sky130_fd_sc_hd__and2_1 _13133_ (.A(net873),
    .B(net982),
    .X(_01210_));
 sky130_fd_sc_hd__and2_1 _13134_ (.A(net870),
    .B(net974),
    .X(_01211_));
 sky130_fd_sc_hd__and2_1 _13135_ (.A(net874),
    .B(net942),
    .X(_01212_));
 sky130_fd_sc_hd__and2_1 _13136_ (.A(net874),
    .B(net996),
    .X(_01213_));
 sky130_fd_sc_hd__and2_1 _13137_ (.A(net873),
    .B(net1036),
    .X(_01214_));
 sky130_fd_sc_hd__and2_1 _13138_ (.A(net874),
    .B(net1066),
    .X(_01215_));
 sky130_fd_sc_hd__and2_1 _13139_ (.A(net876),
    .B(net1602),
    .X(_01216_));
 sky130_fd_sc_hd__nor2_1 _13140_ (.A(net882),
    .B(_06065_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _13141_ (.A(net883),
    .B(_06089_),
    .Y(_01218_));
 sky130_fd_sc_hd__and2_2 _13142_ (.A(net862),
    .B(_06112_),
    .X(_01219_));
 sky130_fd_sc_hd__nor2_1 _13143_ (.A(net883),
    .B(_06135_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _13144_ (.A(net883),
    .B(_06159_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _13145_ (.A(net883),
    .B(_06183_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _13146_ (.A(net883),
    .B(_06207_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_1 _13147_ (.A(net883),
    .B(_06231_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor2_2 _13148_ (.A(net888),
    .B(_06255_),
    .Y(_01225_));
 sky130_fd_sc_hd__nor2_1 _13149_ (.A(net884),
    .B(_06279_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _13150_ (.A(net888),
    .B(_06303_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_1 _13151_ (.A(net884),
    .B(_06327_),
    .Y(_01228_));
 sky130_fd_sc_hd__nor2_1 _13152_ (.A(net884),
    .B(_06351_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_1 _13153_ (.A(net884),
    .B(_06375_),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _13154_ (.A(net884),
    .B(_06399_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_1 _13155_ (.A(net884),
    .B(_06423_),
    .Y(_01232_));
 sky130_fd_sc_hd__nor2_1 _13156_ (.A(net884),
    .B(_06447_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _13157_ (.A(net884),
    .B(_06471_),
    .Y(_01234_));
 sky130_fd_sc_hd__nor2_1 _13158_ (.A(net884),
    .B(_06495_),
    .Y(_01235_));
 sky130_fd_sc_hd__nor2_1 _13159_ (.A(net884),
    .B(_06519_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _13160_ (.A(net884),
    .B(_06543_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _13161_ (.A(net884),
    .B(_06567_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor2_1 _13162_ (.A(net889),
    .B(_06591_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _13163_ (.A(net889),
    .B(_06615_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_1 _13164_ (.A(net889),
    .B(_06639_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_2 _13165_ (.A(net889),
    .B(_06663_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _13166_ (.A(net887),
    .B(net3661),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _13167_ (.A(net887),
    .B(_06711_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _13168_ (.A(net887),
    .B(_06735_),
    .Y(_01245_));
 sky130_fd_sc_hd__nor2_1 _13169_ (.A(net885),
    .B(_06759_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _13170_ (.A(net885),
    .B(_06783_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _13171_ (.A(net885),
    .B(_06807_),
    .Y(_01248_));
 sky130_fd_sc_hd__and2_1 _13172_ (.A(net846),
    .B(_05989_),
    .X(_01249_));
 sky130_fd_sc_hd__and2_1 _13173_ (.A(net849),
    .B(_06017_),
    .X(_01250_));
 sky130_fd_sc_hd__and2_1 _13174_ (.A(net849),
    .B(_02099_),
    .X(_01251_));
 sky130_fd_sc_hd__and2_1 _13175_ (.A(net850),
    .B(_02163_),
    .X(_01252_));
 sky130_fd_sc_hd__and2_1 _13176_ (.A(net850),
    .B(_02217_),
    .X(_01253_));
 sky130_fd_sc_hd__and2_1 _13177_ (.A(net847),
    .B(_02284_),
    .X(_01254_));
 sky130_fd_sc_hd__and2_1 _13178_ (.A(net846),
    .B(_02347_),
    .X(_01255_));
 sky130_fd_sc_hd__and2_1 _13179_ (.A(net847),
    .B(_02418_),
    .X(_01256_));
 sky130_fd_sc_hd__and2_1 _13180_ (.A(net849),
    .B(_02496_),
    .X(_01257_));
 sky130_fd_sc_hd__and2_1 _13181_ (.A(net849),
    .B(_02584_),
    .X(_01258_));
 sky130_fd_sc_hd__and2_1 _13182_ (.A(net849),
    .B(_02674_),
    .X(_01259_));
 sky130_fd_sc_hd__and2_1 _13183_ (.A(net847),
    .B(_02774_),
    .X(_01260_));
 sky130_fd_sc_hd__and2_1 _13184_ (.A(net848),
    .B(_02874_),
    .X(_01261_));
 sky130_fd_sc_hd__and2_1 _13185_ (.A(net848),
    .B(_02977_),
    .X(_01262_));
 sky130_fd_sc_hd__and2_1 _13186_ (.A(net849),
    .B(_03087_),
    .X(_01263_));
 sky130_fd_sc_hd__and2_1 _13187_ (.A(net848),
    .B(_03198_),
    .X(_01264_));
 sky130_fd_sc_hd__and2_1 _13188_ (.A(net863),
    .B(_03317_),
    .X(_01265_));
 sky130_fd_sc_hd__and2_1 _13189_ (.A(net848),
    .B(_03445_),
    .X(_01266_));
 sky130_fd_sc_hd__and2_1 _13190_ (.A(net864),
    .B(_03578_),
    .X(_01267_));
 sky130_fd_sc_hd__and2_1 _13191_ (.A(net864),
    .B(_03719_),
    .X(_01268_));
 sky130_fd_sc_hd__and2_1 _13192_ (.A(net863),
    .B(_03851_),
    .X(_01269_));
 sky130_fd_sc_hd__and2_1 _13193_ (.A(net864),
    .B(_04003_),
    .X(_01270_));
 sky130_fd_sc_hd__and2_1 _13194_ (.A(net865),
    .B(_04151_),
    .X(_01271_));
 sky130_fd_sc_hd__and2_1 _13195_ (.A(net864),
    .B(_04301_),
    .X(_01272_));
 sky130_fd_sc_hd__and2_1 _13196_ (.A(net864),
    .B(_04452_),
    .X(_01273_));
 sky130_fd_sc_hd__and2_1 _13197_ (.A(net865),
    .B(_04627_),
    .X(_01274_));
 sky130_fd_sc_hd__and2_1 _13198_ (.A(net865),
    .B(_04789_),
    .X(_01275_));
 sky130_fd_sc_hd__and2_1 _13199_ (.A(net865),
    .B(_04968_),
    .X(_01276_));
 sky130_fd_sc_hd__and2_1 _13200_ (.A(net879),
    .B(_05139_),
    .X(_01277_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(net865),
    .B(_05328_),
    .X(_01278_));
 sky130_fd_sc_hd__and2_1 _13202_ (.A(net865),
    .B(_05509_),
    .X(_01279_));
 sky130_fd_sc_hd__and2_1 _13203_ (.A(net865),
    .B(_05700_),
    .X(_01280_));
 sky130_fd_sc_hd__nor2_4 _13204_ (.A(_01823_),
    .B(_02024_),
    .Y(_06809_));
 sky130_fd_sc_hd__mux2_1 _13205_ (.A0(net1934),
    .A1(net718),
    .S(net421),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _13206_ (.A0(net3122),
    .A1(net717),
    .S(net421),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _13207_ (.A0(net3006),
    .A1(net714),
    .S(net421),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(net1830),
    .A1(net712),
    .S(net421),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _13209_ (.A0(net1992),
    .A1(net710),
    .S(net421),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _13210_ (.A0(net2368),
    .A1(net708),
    .S(net421),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _13211_ (.A0(net1916),
    .A1(net707),
    .S(net421),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(net2948),
    .A1(net704),
    .S(net421),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(net1422),
    .A1(net703),
    .S(net421),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _13214_ (.A0(net1784),
    .A1(net700),
    .S(net421),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _13215_ (.A0(net1926),
    .A1(net699),
    .S(net421),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _13216_ (.A0(net1876),
    .A1(net697),
    .S(net421),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(net2992),
    .A1(net694),
    .S(net421),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _13218_ (.A0(net1822),
    .A1(net693),
    .S(net421),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(net2436),
    .A1(net690),
    .S(net421),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _13220_ (.A0(net2154),
    .A1(net688),
    .S(net421),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(net1838),
    .A1(net686),
    .S(net422),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _13222_ (.A0(net1242),
    .A1(net684),
    .S(net422),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(net1584),
    .A1(net682),
    .S(net422),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _13224_ (.A0(net1912),
    .A1(net680),
    .S(net422),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(net1202),
    .A1(net677),
    .S(net422),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(net2066),
    .A1(net675),
    .S(net422),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(net1732),
    .A1(net673),
    .S(net422),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _13228_ (.A0(net2652),
    .A1(net671),
    .S(net422),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _13229_ (.A0(net1636),
    .A1(net669),
    .S(net422),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(net1288),
    .A1(\dpath.RF.wdata[25] ),
    .S(net422),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(net1418),
    .A1(net665),
    .S(net422),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(net1448),
    .A1(net663),
    .S(net422),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _13233_ (.A0(net1306),
    .A1(net661),
    .S(net422),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _13234_ (.A0(net1648),
    .A1(net658),
    .S(net422),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _13235_ (.A0(net1346),
    .A1(net657),
    .S(net422),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _13236_ (.A0(net1430),
    .A1(net654),
    .S(net422),
    .X(_01312_));
 sky130_fd_sc_hd__nor2_1 _13237_ (.A(\ctrl.d2c_inst[25] ),
    .B(\ctrl.d2c_inst[24] ),
    .Y(_06810_));
 sky130_fd_sc_hd__and4_1 _13238_ (.A(\ctrl.d2c_inst[31] ),
    .B(\ctrl.d2c_inst[30] ),
    .C(\ctrl.d2c_inst[29] ),
    .D(\ctrl.d2c_inst[28] ),
    .X(_06811_));
 sky130_fd_sc_hd__and4_1 _13239_ (.A(\ctrl.d2c_inst[27] ),
    .B(\ctrl.d2c_inst[26] ),
    .C(_06810_),
    .D(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__and4_4 _13240_ (.A(_01750_),
    .B(\ctrl.d2c_inst[22] ),
    .C(_06026_),
    .D(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__and4_4 _13241_ (.A(net3393),
    .B(net3490),
    .C(_06025_),
    .D(_06812_),
    .X(_06814_));
 sky130_fd_sc_hd__nor2_1 _13242_ (.A(net3724),
    .B(net3722),
    .Y(_06815_));
 sky130_fd_sc_hd__a22o_1 _13243_ (.A1(net129),
    .A2(net3724),
    .B1(net3722),
    .B2(net97),
    .X(_06816_));
 sky130_fd_sc_hd__a21oi_1 _13244_ (.A1(net65),
    .A2(net3719),
    .B1(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__nor2_1 _13245_ (.A(net892),
    .B(_06817_),
    .Y(_01313_));
 sky130_fd_sc_hd__a22o_1 _13246_ (.A1(net140),
    .A2(net3724),
    .B1(net3722),
    .B2(net108),
    .X(_06818_));
 sky130_fd_sc_hd__a21oi_1 _13247_ (.A1(net76),
    .A2(net3719),
    .B1(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__nor2_1 _13248_ (.A(net892),
    .B(_06819_),
    .Y(_01314_));
 sky130_fd_sc_hd__a22o_1 _13249_ (.A1(net151),
    .A2(net3724),
    .B1(net3722),
    .B2(net119),
    .X(_06820_));
 sky130_fd_sc_hd__a21oi_1 _13250_ (.A1(net87),
    .A2(net3719),
    .B1(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__nor2_1 _13251_ (.A(net892),
    .B(_06821_),
    .Y(_01315_));
 sky130_fd_sc_hd__a22o_1 _13252_ (.A1(net154),
    .A2(net3724),
    .B1(net3722),
    .B2(net122),
    .X(_06822_));
 sky130_fd_sc_hd__a21oi_1 _13253_ (.A1(net90),
    .A2(net3719),
    .B1(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__nor2_1 _13254_ (.A(net892),
    .B(_06823_),
    .Y(_01316_));
 sky130_fd_sc_hd__a22o_1 _13255_ (.A1(net155),
    .A2(net3724),
    .B1(net3722),
    .B2(net123),
    .X(_06824_));
 sky130_fd_sc_hd__a21oi_1 _13256_ (.A1(net91),
    .A2(net3719),
    .B1(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__nor2_1 _13257_ (.A(net892),
    .B(_06825_),
    .Y(_01317_));
 sky130_fd_sc_hd__a22o_1 _13258_ (.A1(net156),
    .A2(net3724),
    .B1(net3722),
    .B2(net124),
    .X(_06826_));
 sky130_fd_sc_hd__a21oi_1 _13259_ (.A1(net92),
    .A2(net3719),
    .B1(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__nor2_1 _13260_ (.A(net892),
    .B(_06827_),
    .Y(_01318_));
 sky130_fd_sc_hd__a22o_1 _13261_ (.A1(net157),
    .A2(net3724),
    .B1(net3722),
    .B2(net125),
    .X(_06828_));
 sky130_fd_sc_hd__a21oi_1 _13262_ (.A1(net93),
    .A2(net3719),
    .B1(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__nor2_1 _13263_ (.A(net892),
    .B(_06829_),
    .Y(_01319_));
 sky130_fd_sc_hd__a22o_1 _13264_ (.A1(net158),
    .A2(net3724),
    .B1(net3722),
    .B2(net126),
    .X(_06830_));
 sky130_fd_sc_hd__a21oi_1 _13265_ (.A1(net94),
    .A2(net3719),
    .B1(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__nor2_1 _13266_ (.A(net892),
    .B(_06831_),
    .Y(_01320_));
 sky130_fd_sc_hd__a22o_1 _13267_ (.A1(net159),
    .A2(net3724),
    .B1(net3722),
    .B2(net127),
    .X(_06832_));
 sky130_fd_sc_hd__a21oi_1 _13268_ (.A1(net95),
    .A2(net3719),
    .B1(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__nor2_1 _13269_ (.A(net892),
    .B(_06833_),
    .Y(_01321_));
 sky130_fd_sc_hd__a22o_1 _13270_ (.A1(net160),
    .A2(net3724),
    .B1(net3722),
    .B2(net128),
    .X(_06834_));
 sky130_fd_sc_hd__a21oi_1 _13271_ (.A1(net96),
    .A2(net3719),
    .B1(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__nor2_1 _13272_ (.A(net892),
    .B(_06835_),
    .Y(_01322_));
 sky130_fd_sc_hd__a22o_1 _13273_ (.A1(net130),
    .A2(net3724),
    .B1(net3722),
    .B2(net98),
    .X(_06836_));
 sky130_fd_sc_hd__a21oi_1 _13274_ (.A1(net66),
    .A2(net3719),
    .B1(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__nor2_1 _13275_ (.A(net892),
    .B(_06837_),
    .Y(_01323_));
 sky130_fd_sc_hd__a22o_1 _13276_ (.A1(net131),
    .A2(net3724),
    .B1(net3722),
    .B2(net99),
    .X(_06838_));
 sky130_fd_sc_hd__a21oi_1 _13277_ (.A1(net67),
    .A2(net3719),
    .B1(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__nor2_1 _13278_ (.A(net892),
    .B(_06839_),
    .Y(_01324_));
 sky130_fd_sc_hd__a22o_1 _13279_ (.A1(net132),
    .A2(net3724),
    .B1(net3722),
    .B2(net100),
    .X(_06840_));
 sky130_fd_sc_hd__a21oi_1 _13280_ (.A1(net68),
    .A2(net3719),
    .B1(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__nor2_1 _13281_ (.A(net892),
    .B(_06841_),
    .Y(_01325_));
 sky130_fd_sc_hd__a22o_1 _13282_ (.A1(net133),
    .A2(net3724),
    .B1(net3722),
    .B2(net101),
    .X(_06842_));
 sky130_fd_sc_hd__a21oi_1 _13283_ (.A1(net69),
    .A2(net3719),
    .B1(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__nor2_1 _13284_ (.A(net892),
    .B(_06843_),
    .Y(_01326_));
 sky130_fd_sc_hd__a22o_1 _13285_ (.A1(net134),
    .A2(net3724),
    .B1(net3722),
    .B2(net102),
    .X(_06844_));
 sky130_fd_sc_hd__a21oi_1 _13286_ (.A1(net70),
    .A2(net3719),
    .B1(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__nor2_1 _13287_ (.A(net892),
    .B(_06845_),
    .Y(_01327_));
 sky130_fd_sc_hd__a22o_1 _13288_ (.A1(net135),
    .A2(net3723),
    .B1(net3721),
    .B2(net103),
    .X(_06846_));
 sky130_fd_sc_hd__a21oi_1 _13289_ (.A1(net71),
    .A2(net3719),
    .B1(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__nor2_1 _13290_ (.A(net893),
    .B(_06847_),
    .Y(_01328_));
 sky130_fd_sc_hd__a22o_1 _13291_ (.A1(net136),
    .A2(net3723),
    .B1(net3721),
    .B2(net104),
    .X(_06848_));
 sky130_fd_sc_hd__a21oi_1 _13292_ (.A1(net72),
    .A2(net3720),
    .B1(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__nor2_1 _13293_ (.A(net893),
    .B(_06849_),
    .Y(_01329_));
 sky130_fd_sc_hd__a22o_1 _13294_ (.A1(net137),
    .A2(net3723),
    .B1(net3721),
    .B2(net105),
    .X(_06850_));
 sky130_fd_sc_hd__a21oi_1 _13295_ (.A1(net73),
    .A2(net3720),
    .B1(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__nor2_1 _13296_ (.A(net893),
    .B(_06851_),
    .Y(_01330_));
 sky130_fd_sc_hd__a22o_1 _13297_ (.A1(net138),
    .A2(net3723),
    .B1(net3721),
    .B2(net106),
    .X(_06852_));
 sky130_fd_sc_hd__a21oi_1 _13298_ (.A1(net74),
    .A2(net3720),
    .B1(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__nor2_1 _13299_ (.A(net893),
    .B(_06853_),
    .Y(_01331_));
 sky130_fd_sc_hd__a22o_1 _13300_ (.A1(net139),
    .A2(net3723),
    .B1(net3721),
    .B2(net107),
    .X(_06854_));
 sky130_fd_sc_hd__a21oi_1 _13301_ (.A1(net75),
    .A2(net3720),
    .B1(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__nor2_1 _13302_ (.A(net893),
    .B(_06855_),
    .Y(_01332_));
 sky130_fd_sc_hd__a22o_1 _13303_ (.A1(net141),
    .A2(net3723),
    .B1(net3721),
    .B2(net109),
    .X(_06856_));
 sky130_fd_sc_hd__a21oi_1 _13304_ (.A1(net77),
    .A2(net3720),
    .B1(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2_1 _13305_ (.A(net893),
    .B(_06857_),
    .Y(_01333_));
 sky130_fd_sc_hd__a22o_1 _13306_ (.A1(net142),
    .A2(net3723),
    .B1(net3721),
    .B2(net110),
    .X(_06858_));
 sky130_fd_sc_hd__a21oi_1 _13307_ (.A1(net78),
    .A2(net3720),
    .B1(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__nor2_1 _13308_ (.A(net893),
    .B(_06859_),
    .Y(_01334_));
 sky130_fd_sc_hd__a22o_1 _13309_ (.A1(net143),
    .A2(net3723),
    .B1(net3721),
    .B2(net111),
    .X(_06860_));
 sky130_fd_sc_hd__a21oi_1 _13310_ (.A1(net79),
    .A2(net3720),
    .B1(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__nor2_1 _13311_ (.A(net893),
    .B(_06861_),
    .Y(_01335_));
 sky130_fd_sc_hd__a22o_1 _13312_ (.A1(net144),
    .A2(net3723),
    .B1(net3721),
    .B2(net112),
    .X(_06862_));
 sky130_fd_sc_hd__a21oi_1 _13313_ (.A1(net80),
    .A2(net3720),
    .B1(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__nor2_1 _13314_ (.A(net893),
    .B(_06863_),
    .Y(_01336_));
 sky130_fd_sc_hd__a22o_1 _13315_ (.A1(net145),
    .A2(net3723),
    .B1(net3721),
    .B2(net113),
    .X(_06864_));
 sky130_fd_sc_hd__a21oi_1 _13316_ (.A1(net81),
    .A2(net3720),
    .B1(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__nor2_1 _13317_ (.A(net893),
    .B(_06865_),
    .Y(_01337_));
 sky130_fd_sc_hd__a22o_1 _13318_ (.A1(net146),
    .A2(net3723),
    .B1(net3721),
    .B2(net114),
    .X(_06866_));
 sky130_fd_sc_hd__a21oi_1 _13319_ (.A1(net82),
    .A2(net3720),
    .B1(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__nor2_1 _13320_ (.A(net894),
    .B(_06867_),
    .Y(_01338_));
 sky130_fd_sc_hd__a22o_1 _13321_ (.A1(net147),
    .A2(net3723),
    .B1(net3721),
    .B2(net115),
    .X(_06868_));
 sky130_fd_sc_hd__a21oi_1 _13322_ (.A1(net83),
    .A2(net3720),
    .B1(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__nor2_1 _13323_ (.A(net894),
    .B(_06869_),
    .Y(_01339_));
 sky130_fd_sc_hd__a22o_1 _13324_ (.A1(net148),
    .A2(net3723),
    .B1(net3721),
    .B2(net116),
    .X(_06870_));
 sky130_fd_sc_hd__a21oi_1 _13325_ (.A1(net84),
    .A2(net3720),
    .B1(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__nor2_1 _13326_ (.A(net894),
    .B(_06871_),
    .Y(_01340_));
 sky130_fd_sc_hd__a22o_1 _13327_ (.A1(net149),
    .A2(net3723),
    .B1(net3721),
    .B2(net117),
    .X(_06872_));
 sky130_fd_sc_hd__a21oi_1 _13328_ (.A1(net85),
    .A2(net3720),
    .B1(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nor2_1 _13329_ (.A(net894),
    .B(_06873_),
    .Y(_01341_));
 sky130_fd_sc_hd__a22o_1 _13330_ (.A1(net150),
    .A2(net3723),
    .B1(net3721),
    .B2(net118),
    .X(_06874_));
 sky130_fd_sc_hd__a21oi_1 _13331_ (.A1(net86),
    .A2(net3720),
    .B1(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__nor2_1 _13332_ (.A(net894),
    .B(_06875_),
    .Y(_01342_));
 sky130_fd_sc_hd__a22o_1 _13333_ (.A1(net152),
    .A2(_06813_),
    .B1(_06814_),
    .B2(net120),
    .X(_06876_));
 sky130_fd_sc_hd__a21oi_1 _13334_ (.A1(net88),
    .A2(net3720),
    .B1(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__nor2_1 _13335_ (.A(net894),
    .B(_06877_),
    .Y(_01343_));
 sky130_fd_sc_hd__a22o_1 _13336_ (.A1(net153),
    .A2(net3723),
    .B1(net3721),
    .B2(net121),
    .X(_06878_));
 sky130_fd_sc_hd__a21oi_1 _13337_ (.A1(net89),
    .A2(net3720),
    .B1(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nor2_1 _13338_ (.A(net894),
    .B(_06879_),
    .Y(_01344_));
 sky130_fd_sc_hd__a21oi_1 _13339_ (.A1(_02125_),
    .A2(_02128_),
    .B1(net3249),
    .Y(_06880_));
 sky130_fd_sc_hd__or2_1 _13340_ (.A(_02129_),
    .B(net3250),
    .X(_06881_));
 sky130_fd_sc_hd__nor2_1 _13341_ (.A(net880),
    .B(net3251),
    .Y(_01345_));
 sky130_fd_sc_hd__xor2_1 _13342_ (.A(_02129_),
    .B(_02131_),
    .X(_06882_));
 sky130_fd_sc_hd__nor2_1 _13343_ (.A(net880),
    .B(_06882_),
    .Y(_01346_));
 sky130_fd_sc_hd__nor2_1 _13344_ (.A(net880),
    .B(_02137_),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2_1 _13345_ (.A(net880),
    .B(_02191_),
    .Y(_01348_));
 sky130_fd_sc_hd__nor2_1 _13346_ (.A(net881),
    .B(_02254_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_1 _13347_ (.A(net881),
    .B(_02322_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_1 _13348_ (.A(net881),
    .B(_02393_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _13349_ (.A(net881),
    .B(_02466_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _13350_ (.A(net881),
    .B(_02557_),
    .Y(_01353_));
 sky130_fd_sc_hd__nor2_1 _13351_ (.A(net881),
    .B(_02646_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_1 _13352_ (.A(net881),
    .B(_02746_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _13353_ (.A(net881),
    .B(_02849_),
    .Y(_01356_));
 sky130_fd_sc_hd__nor2_1 _13354_ (.A(net881),
    .B(_02952_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _13355_ (.A(net881),
    .B(_03059_),
    .Y(_01358_));
 sky130_fd_sc_hd__nor2_1 _13356_ (.A(net881),
    .B(_03173_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _13357_ (.A(net881),
    .B(_03289_),
    .Y(_01360_));
 sky130_fd_sc_hd__nor2_1 _13358_ (.A(net881),
    .B(_03420_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _13359_ (.A(net881),
    .B(_03550_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_1 _13360_ (.A(net881),
    .B(_03691_),
    .Y(_01363_));
 sky130_fd_sc_hd__nor2_1 _13361_ (.A(net880),
    .B(_03827_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _13362_ (.A(net880),
    .B(_03976_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _13363_ (.A(net880),
    .B(_04118_),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_1 _13364_ (.A(net880),
    .B(_04129_),
    .Y(_01367_));
 sky130_fd_sc_hd__nor2_1 _13365_ (.A(net880),
    .B(_04425_),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _13366_ (.A(net880),
    .B(_04601_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_1 _13367_ (.A(net880),
    .B(_04763_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _13368_ (.A(net880),
    .B(_04941_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _13369_ (.A(net880),
    .B(_05114_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _13370_ (.A(net882),
    .B(_05302_),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_1 _13371_ (.A(net882),
    .B(_05483_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _13372_ (.A(net882),
    .B(_05672_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor3_1 _13373_ (.A(net882),
    .B(_05833_),
    .C(_05834_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _13374_ (.A(net883),
    .B(_05987_),
    .Y(_01377_));
 sky130_fd_sc_hd__and2_1 _13375_ (.A(net850),
    .B(_06022_),
    .X(_01378_));
 sky130_fd_sc_hd__and2_1 _13376_ (.A(net850),
    .B(_02114_),
    .X(_01379_));
 sky130_fd_sc_hd__and2_1 _13377_ (.A(net850),
    .B(_02183_),
    .X(_01380_));
 sky130_fd_sc_hd__and2_1 _13378_ (.A(net850),
    .B(_02246_),
    .X(_01381_));
 sky130_fd_sc_hd__and2_1 _13379_ (.A(net847),
    .B(_02316_),
    .X(_01382_));
 sky130_fd_sc_hd__nor2_1 _13380_ (.A(net883),
    .B(_02386_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _13381_ (.A(net883),
    .B(_02458_),
    .Y(_01384_));
 sky130_fd_sc_hd__and2_1 _13382_ (.A(net847),
    .B(_02551_),
    .X(_01385_));
 sky130_fd_sc_hd__and2_1 _13383_ (.A(net847),
    .B(_02640_),
    .X(_01386_));
 sky130_fd_sc_hd__nor2_1 _13384_ (.A(net884),
    .B(_02739_),
    .Y(_01387_));
 sky130_fd_sc_hd__and2_1 _13385_ (.A(net847),
    .B(_02840_),
    .X(_01388_));
 sky130_fd_sc_hd__and2_1 _13386_ (.A(net847),
    .B(_02944_),
    .X(_01389_));
 sky130_fd_sc_hd__and2_1 _13387_ (.A(net848),
    .B(_03052_),
    .X(_01390_));
 sky130_fd_sc_hd__and2_1 _13388_ (.A(net848),
    .B(_03166_),
    .X(_01391_));
 sky130_fd_sc_hd__nor2_1 _13389_ (.A(net884),
    .B(_03281_),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _13390_ (.A(net889),
    .B(_03410_),
    .Y(_01393_));
 sky130_fd_sc_hd__and2_1 _13391_ (.A(net848),
    .B(net3673),
    .X(_01394_));
 sky130_fd_sc_hd__and2_1 _13392_ (.A(net863),
    .B(_03684_),
    .X(_01395_));
 sky130_fd_sc_hd__and2_1 _13393_ (.A(net848),
    .B(_03820_),
    .X(_01396_));
 sky130_fd_sc_hd__and2_1 _13394_ (.A(net864),
    .B(_03968_),
    .X(_01397_));
 sky130_fd_sc_hd__and2_1 _13395_ (.A(net863),
    .B(_04113_),
    .X(_01398_));
 sky130_fd_sc_hd__and2_1 _13396_ (.A(net863),
    .B(_04275_),
    .X(_01399_));
 sky130_fd_sc_hd__and2_1 _13397_ (.A(net864),
    .B(_04421_),
    .X(_01400_));
 sky130_fd_sc_hd__and2_2 _13398_ (.A(net879),
    .B(_04593_),
    .X(_01401_));
 sky130_fd_sc_hd__and2_1 _13399_ (.A(net865),
    .B(net3692),
    .X(_01402_));
 sky130_fd_sc_hd__and2_1 _13400_ (.A(net849),
    .B(net3602),
    .X(_01403_));
 sky130_fd_sc_hd__and2_1 _13401_ (.A(net865),
    .B(net3647),
    .X(_01404_));
 sky130_fd_sc_hd__and2_1 _13402_ (.A(net879),
    .B(net3610),
    .X(_01405_));
 sky130_fd_sc_hd__and2_1 _13403_ (.A(net865),
    .B(net3675),
    .X(_01406_));
 sky130_fd_sc_hd__and2_1 _13404_ (.A(net865),
    .B(net3337),
    .X(_01407_));
 sky130_fd_sc_hd__and2_1 _13405_ (.A(net879),
    .B(net3680),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _13406_ (.A(net475),
    .B(net3311),
    .Y(_06883_));
 sky130_fd_sc_hd__o211a_1 _13407_ (.A1(net3249),
    .A2(net475),
    .B1(_06883_),
    .C1(net852),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _13408_ (.A0(net3233),
    .A1(_06024_),
    .S(net475),
    .X(_06884_));
 sky130_fd_sc_hd__and2_1 _13409_ (.A(net852),
    .B(_06884_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _13410_ (.A0(net3518),
    .A1(_02118_),
    .S(net475),
    .X(_06885_));
 sky130_fd_sc_hd__and2_1 _13411_ (.A(net858),
    .B(_06885_),
    .X(_01411_));
 sky130_fd_sc_hd__nand2_1 _13412_ (.A(net474),
    .B(net3273),
    .Y(_06886_));
 sky130_fd_sc_hd__o211a_1 _13413_ (.A1(net3231),
    .A2(net474),
    .B1(_06886_),
    .C1(net846),
    .X(_01412_));
 sky130_fd_sc_hd__nand2_1 _13414_ (.A(net476),
    .B(net3269),
    .Y(_06887_));
 sky130_fd_sc_hd__o211a_1 _13415_ (.A1(net3238),
    .A2(net476),
    .B1(_06887_),
    .C1(net846),
    .X(_01413_));
 sky130_fd_sc_hd__nand2_1 _13416_ (.A(net476),
    .B(_02317_),
    .Y(_06888_));
 sky130_fd_sc_hd__o211a_1 _13417_ (.A1(net1338),
    .A2(net476),
    .B1(_06888_),
    .C1(net846),
    .X(_01414_));
 sky130_fd_sc_hd__nand2_1 _13418_ (.A(net476),
    .B(net3412),
    .Y(_06889_));
 sky130_fd_sc_hd__o211a_1 _13419_ (.A1(net3297),
    .A2(net476),
    .B1(_06889_),
    .C1(net846),
    .X(_01415_));
 sky130_fd_sc_hd__nand2_1 _13420_ (.A(net473),
    .B(net3400),
    .Y(_06890_));
 sky130_fd_sc_hd__o211a_1 _13421_ (.A1(net3277),
    .A2(net473),
    .B1(_06890_),
    .C1(net846),
    .X(_01416_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(net474),
    .B(net3417),
    .Y(_06891_));
 sky130_fd_sc_hd__o211a_1 _13423_ (.A1(net3286),
    .A2(net474),
    .B1(_06891_),
    .C1(net846),
    .X(_01417_));
 sky130_fd_sc_hd__nand2_1 _13424_ (.A(net473),
    .B(_02641_),
    .Y(_06892_));
 sky130_fd_sc_hd__o211a_1 _13425_ (.A1(net3228),
    .A2(net474),
    .B1(_06892_),
    .C1(net843),
    .X(_01418_));
 sky130_fd_sc_hd__nand2_1 _13426_ (.A(net473),
    .B(net3485),
    .Y(_06893_));
 sky130_fd_sc_hd__o211a_1 _13427_ (.A1(net3274),
    .A2(net473),
    .B1(_06893_),
    .C1(net843),
    .X(_01419_));
 sky130_fd_sc_hd__nand2_1 _13428_ (.A(net473),
    .B(_02841_),
    .Y(_06894_));
 sky130_fd_sc_hd__o211a_1 _13429_ (.A1(net3358),
    .A2(net473),
    .B1(_06894_),
    .C1(net843),
    .X(_01420_));
 sky130_fd_sc_hd__nand2_1 _13430_ (.A(net473),
    .B(_02945_),
    .Y(_06895_));
 sky130_fd_sc_hd__o211a_1 _13431_ (.A1(net3301),
    .A2(net473),
    .B1(_06895_),
    .C1(net843),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(net3295),
    .A1(_03053_),
    .S(net473),
    .X(_06896_));
 sky130_fd_sc_hd__and2_1 _13433_ (.A(net843),
    .B(_06896_),
    .X(_01422_));
 sky130_fd_sc_hd__nand2_1 _13434_ (.A(net473),
    .B(_03167_),
    .Y(_06897_));
 sky130_fd_sc_hd__o211a_2 _13435_ (.A1(net3291),
    .A2(net473),
    .B1(_06897_),
    .C1(net843),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_2 _13436_ (.A0(net3241),
    .A1(_03283_),
    .S(net473),
    .X(_06898_));
 sky130_fd_sc_hd__and2_1 _13437_ (.A(net862),
    .B(_06898_),
    .X(_01424_));
 sky130_fd_sc_hd__nand2_1 _13438_ (.A(net473),
    .B(net3454),
    .Y(_06899_));
 sky130_fd_sc_hd__o211a_1 _13439_ (.A1(net3265),
    .A2(net473),
    .B1(_06899_),
    .C1(net843),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_2 _13440_ (.A0(net3221),
    .A1(_03544_),
    .S(net473),
    .X(_06900_));
 sky130_fd_sc_hd__and2_1 _13441_ (.A(net858),
    .B(_06900_),
    .X(_01426_));
 sky130_fd_sc_hd__nand2_1 _13442_ (.A(net474),
    .B(_03685_),
    .Y(_06901_));
 sky130_fd_sc_hd__o211a_1 _13443_ (.A1(net3325),
    .A2(net474),
    .B1(_06901_),
    .C1(net843),
    .X(_01427_));
 sky130_fd_sc_hd__nand2_1 _13444_ (.A(net474),
    .B(_03821_),
    .Y(_06902_));
 sky130_fd_sc_hd__o211a_1 _13445_ (.A1(net3323),
    .A2(net474),
    .B1(_06902_),
    .C1(net844),
    .X(_01428_));
 sky130_fd_sc_hd__nand2_1 _13446_ (.A(net474),
    .B(_03969_),
    .Y(_01673_));
 sky130_fd_sc_hd__o211a_1 _13447_ (.A1(net3462),
    .A2(net474),
    .B1(_01673_),
    .C1(net843),
    .X(_01429_));
 sky130_fd_sc_hd__nand2_1 _13448_ (.A(net474),
    .B(_04114_),
    .Y(_01674_));
 sky130_fd_sc_hd__o211a_1 _13449_ (.A1(net3455),
    .A2(net474),
    .B1(_01674_),
    .C1(net843),
    .X(_01430_));
 sky130_fd_sc_hd__nand2_1 _13450_ (.A(net474),
    .B(_04276_),
    .Y(_01675_));
 sky130_fd_sc_hd__o211a_1 _13451_ (.A1(net3466),
    .A2(net475),
    .B1(_01675_),
    .C1(net852),
    .X(_01431_));
 sky130_fd_sc_hd__nand2_1 _13452_ (.A(net475),
    .B(_04422_),
    .Y(_01676_));
 sky130_fd_sc_hd__o211a_1 _13453_ (.A1(net3468),
    .A2(net475),
    .B1(_01676_),
    .C1(net851),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(net3542),
    .A1(_04594_),
    .S(net475),
    .X(_01677_));
 sky130_fd_sc_hd__and2_1 _13455_ (.A(net862),
    .B(_01677_),
    .X(_01433_));
 sky130_fd_sc_hd__nand2_1 _13456_ (.A(net475),
    .B(_04760_),
    .Y(_01678_));
 sky130_fd_sc_hd__o211a_1 _13457_ (.A1(net3522),
    .A2(net476),
    .B1(_01678_),
    .C1(net858),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _13458_ (.A0(net3509),
    .A1(_04934_),
    .S(net476),
    .X(_01679_));
 sky130_fd_sc_hd__and2_1 _13459_ (.A(net858),
    .B(_01679_),
    .X(_01435_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(net475),
    .B(_05110_),
    .Y(_01680_));
 sky130_fd_sc_hd__o211a_1 _13461_ (.A1(net3339),
    .A2(net475),
    .B1(_01680_),
    .C1(net858),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _13462_ (.A0(net3401),
    .A1(_05293_),
    .S(net475),
    .X(_01681_));
 sky130_fd_sc_hd__and2_1 _13463_ (.A(net857),
    .B(_01681_),
    .X(_01437_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(net476),
    .B(_05477_),
    .Y(_01682_));
 sky130_fd_sc_hd__o211a_1 _13465_ (.A1(net3439),
    .A2(net475),
    .B1(_01682_),
    .C1(net858),
    .X(_01438_));
 sky130_fd_sc_hd__nand2_1 _13466_ (.A(net476),
    .B(_05663_),
    .Y(_01683_));
 sky130_fd_sc_hd__o211a_1 _13467_ (.A1(net3283),
    .A2(net476),
    .B1(_01683_),
    .C1(net858),
    .X(_01439_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(net475),
    .B(_05829_),
    .Y(_01684_));
 sky130_fd_sc_hd__o211a_1 _13469_ (.A1(net3184),
    .A2(net475),
    .B1(_01684_),
    .C1(net858),
    .X(_01440_));
 sky130_fd_sc_hd__and2_1 _13470_ (.A(net876),
    .B(net1140),
    .X(_01441_));
 sky130_fd_sc_hd__and2_1 _13471_ (.A(net879),
    .B(net2620),
    .X(_01442_));
 sky130_fd_sc_hd__and2_1 _13472_ (.A(net849),
    .B(net3170),
    .X(_01443_));
 sky130_fd_sc_hd__and2_2 _13473_ (.A(net849),
    .B(net3194),
    .X(_01444_));
 sky130_fd_sc_hd__and2_2 _13474_ (.A(net849),
    .B(net3230),
    .X(_01445_));
 sky130_fd_sc_hd__and2_1 _13475_ (.A(net849),
    .B(net2092),
    .X(_01446_));
 sky130_fd_sc_hd__and2_2 _13476_ (.A(net849),
    .B(net3210),
    .X(_01447_));
 sky130_fd_sc_hd__and2_1 _13477_ (.A(net850),
    .B(net3178),
    .X(_01448_));
 sky130_fd_sc_hd__and2_1 _13478_ (.A(net871),
    .B(net902),
    .X(_01449_));
 sky130_fd_sc_hd__and2_1 _13479_ (.A(net879),
    .B(net3220),
    .X(_01450_));
 sky130_fd_sc_hd__and2_1 _13480_ (.A(net870),
    .B(net1018),
    .X(_01451_));
 sky130_fd_sc_hd__and2_1 _13481_ (.A(net849),
    .B(net1970),
    .X(_01452_));
 sky130_fd_sc_hd__and2_1 _13482_ (.A(net868),
    .B(net898),
    .X(_01453_));
 sky130_fd_sc_hd__and2_1 _13483_ (.A(net871),
    .B(net1002),
    .X(_01454_));
 sky130_fd_sc_hd__and2_1 _13484_ (.A(net868),
    .B(net992),
    .X(_01455_));
 sky130_fd_sc_hd__and2_1 _13485_ (.A(net870),
    .B(net980),
    .X(_01456_));
 sky130_fd_sc_hd__and2_1 _13486_ (.A(net872),
    .B(net1016),
    .X(_01457_));
 sky130_fd_sc_hd__and2_1 _13487_ (.A(net871),
    .B(net904),
    .X(_01458_));
 sky130_fd_sc_hd__and2_1 _13488_ (.A(net868),
    .B(net984),
    .X(_01459_));
 sky130_fd_sc_hd__and2_1 _13489_ (.A(net869),
    .B(net930),
    .X(_01460_));
 sky130_fd_sc_hd__and2_1 _13490_ (.A(net868),
    .B(net954),
    .X(_01461_));
 sky130_fd_sc_hd__and2_1 _13491_ (.A(net867),
    .B(net948),
    .X(_01462_));
 sky130_fd_sc_hd__and2_1 _13492_ (.A(net870),
    .B(net952),
    .X(_01463_));
 sky130_fd_sc_hd__and2_1 _13493_ (.A(net873),
    .B(net1028),
    .X(_01464_));
 sky130_fd_sc_hd__and2_1 _13494_ (.A(net874),
    .B(net936),
    .X(_01465_));
 sky130_fd_sc_hd__and2_1 _13495_ (.A(net873),
    .B(net918),
    .X(_01466_));
 sky130_fd_sc_hd__and2_1 _13496_ (.A(net874),
    .B(net994),
    .X(_01467_));
 sky130_fd_sc_hd__and2_1 _13497_ (.A(net874),
    .B(net1004),
    .X(_01468_));
 sky130_fd_sc_hd__and2_1 _13498_ (.A(net874),
    .B(net938),
    .X(_01469_));
 sky130_fd_sc_hd__and2_1 _13499_ (.A(net874),
    .B(net3062),
    .X(_01470_));
 sky130_fd_sc_hd__and2_1 _13500_ (.A(net876),
    .B(net1008),
    .X(_01471_));
 sky130_fd_sc_hd__and2_1 _13501_ (.A(net876),
    .B(net900),
    .X(_01472_));
 sky130_fd_sc_hd__nand2_4 _13502_ (.A(_01829_),
    .B(_02023_),
    .Y(_01685_));
 sky130_fd_sc_hd__mux2_1 _13503_ (.A0(net718),
    .A1(net3056),
    .S(net375),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(net717),
    .A1(net2250),
    .S(net375),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(net714),
    .A1(net1938),
    .S(net375),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _13506_ (.A0(net712),
    .A1(net3156),
    .S(net375),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _13507_ (.A0(net711),
    .A1(net2906),
    .S(net375),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(net709),
    .A1(net3016),
    .S(net375),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _13509_ (.A0(net706),
    .A1(net2780),
    .S(net375),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(net704),
    .A1(net2832),
    .S(net375),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(net703),
    .A1(net2312),
    .S(net375),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _13512_ (.A0(net700),
    .A1(net2922),
    .S(net375),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _13513_ (.A0(net698),
    .A1(net3044),
    .S(net375),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(net697),
    .A1(net1600),
    .S(net375),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(net694),
    .A1(net2740),
    .S(net375),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(net693),
    .A1(net3190),
    .S(net375),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _13517_ (.A0(net690),
    .A1(net2178),
    .S(net375),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(net688),
    .A1(net1842),
    .S(net375),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(net686),
    .A1(net2208),
    .S(net376),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(net684),
    .A1(net2404),
    .S(net376),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _13521_ (.A0(net682),
    .A1(net3064),
    .S(net376),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _13522_ (.A0(net680),
    .A1(net2300),
    .S(net376),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _13523_ (.A0(net677),
    .A1(net2506),
    .S(net376),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(net675),
    .A1(net2216),
    .S(net376),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _13525_ (.A0(net673),
    .A1(net1846),
    .S(net376),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(net672),
    .A1(net2626),
    .S(net376),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _13527_ (.A0(net669),
    .A1(net1520),
    .S(net376),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(net667),
    .A1(net2968),
    .S(net376),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _13529_ (.A0(net665),
    .A1(net1344),
    .S(net376),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(net663),
    .A1(net2504),
    .S(net376),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _13531_ (.A0(net661),
    .A1(net1858),
    .S(net376),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(net658),
    .A1(net2040),
    .S(net376),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _13533_ (.A0(net657),
    .A1(net1572),
    .S(net376),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(\dpath.RF.wdata[31] ),
    .A1(net1664),
    .S(net376),
    .X(_01504_));
 sky130_fd_sc_hd__and2_1 _13535_ (.A(net3327),
    .B(net857),
    .X(_01505_));
 sky130_fd_sc_hd__or2_1 _13536_ (.A(net3341),
    .B(net452),
    .X(_01686_));
 sky130_fd_sc_hd__o211a_1 _13537_ (.A1(net3249),
    .A2(net445),
    .B1(_01686_),
    .C1(net851),
    .X(_01506_));
 sky130_fd_sc_hd__or2_1 _13538_ (.A(net239),
    .B(net452),
    .X(_01687_));
 sky130_fd_sc_hd__o211a_1 _13539_ (.A1(net3233),
    .A2(net445),
    .B1(_01687_),
    .C1(net852),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(net250),
    .A1(net3518),
    .S(net451),
    .X(_01688_));
 sky130_fd_sc_hd__and2_1 _13541_ (.A(net843),
    .B(net3519),
    .X(_01508_));
 sky130_fd_sc_hd__or2_1 _13542_ (.A(net253),
    .B(net451),
    .X(_01689_));
 sky130_fd_sc_hd__o211a_1 _13543_ (.A1(net3231),
    .A2(net444),
    .B1(_01689_),
    .C1(net843),
    .X(_01509_));
 sky130_fd_sc_hd__or2_1 _13544_ (.A(net254),
    .B(net450),
    .X(_01690_));
 sky130_fd_sc_hd__o211a_1 _13545_ (.A1(net3238),
    .A2(net442),
    .B1(_01690_),
    .C1(net846),
    .X(_01510_));
 sky130_fd_sc_hd__or2_1 _13546_ (.A(net3280),
    .B(net450),
    .X(_01691_));
 sky130_fd_sc_hd__o211a_1 _13547_ (.A1(net1338),
    .A2(net442),
    .B1(_01691_),
    .C1(net846),
    .X(_01511_));
 sky130_fd_sc_hd__or2_1 _13548_ (.A(net256),
    .B(net450),
    .X(_01692_));
 sky130_fd_sc_hd__o211a_1 _13549_ (.A1(net3297),
    .A2(net442),
    .B1(_01692_),
    .C1(net846),
    .X(_01512_));
 sky130_fd_sc_hd__or2_1 _13550_ (.A(net257),
    .B(net450),
    .X(_01693_));
 sky130_fd_sc_hd__o211a_1 _13551_ (.A1(net3277),
    .A2(net442),
    .B1(_01693_),
    .C1(net843),
    .X(_01513_));
 sky130_fd_sc_hd__or2_1 _13552_ (.A(net258),
    .B(net450),
    .X(_01694_));
 sky130_fd_sc_hd__o211a_1 _13553_ (.A1(net3286),
    .A2(net444),
    .B1(_01694_),
    .C1(net843),
    .X(_01514_));
 sky130_fd_sc_hd__or2_1 _13554_ (.A(net3375),
    .B(net450),
    .X(_01695_));
 sky130_fd_sc_hd__o211a_1 _13555_ (.A1(net3228),
    .A2(net442),
    .B1(_01695_),
    .C1(net845),
    .X(_01515_));
 sky130_fd_sc_hd__or2_1 _13556_ (.A(net229),
    .B(net449),
    .X(_01696_));
 sky130_fd_sc_hd__o211a_1 _13557_ (.A1(net3274),
    .A2(net441),
    .B1(_01696_),
    .C1(net843),
    .X(_01516_));
 sky130_fd_sc_hd__or2_1 _13558_ (.A(net3410),
    .B(net449),
    .X(_01697_));
 sky130_fd_sc_hd__o211a_1 _13559_ (.A1(net3358),
    .A2(net441),
    .B1(_01697_),
    .C1(net845),
    .X(_01517_));
 sky130_fd_sc_hd__or2_1 _13560_ (.A(net231),
    .B(net449),
    .X(_01698_));
 sky130_fd_sc_hd__o211a_1 _13561_ (.A1(net3301),
    .A2(net441),
    .B1(_01698_),
    .C1(net845),
    .X(_01518_));
 sky130_fd_sc_hd__or2_1 _13562_ (.A(net232),
    .B(net449),
    .X(_01699_));
 sky130_fd_sc_hd__o211a_1 _13563_ (.A1(net3295),
    .A2(net441),
    .B1(_01699_),
    .C1(net845),
    .X(_01519_));
 sky130_fd_sc_hd__or2_1 _13564_ (.A(net233),
    .B(net449),
    .X(_01700_));
 sky130_fd_sc_hd__o211a_1 _13565_ (.A1(net3291),
    .A2(net441),
    .B1(_01700_),
    .C1(net845),
    .X(_01520_));
 sky130_fd_sc_hd__or2_1 _13566_ (.A(net234),
    .B(net449),
    .X(_01701_));
 sky130_fd_sc_hd__o211a_1 _13567_ (.A1(net3241),
    .A2(net441),
    .B1(_01701_),
    .C1(net844),
    .X(_01521_));
 sky130_fd_sc_hd__or2_1 _13568_ (.A(net235),
    .B(net449),
    .X(_01702_));
 sky130_fd_sc_hd__o211a_1 _13569_ (.A1(net3265),
    .A2(net442),
    .B1(_01702_),
    .C1(net844),
    .X(_01522_));
 sky130_fd_sc_hd__or2_1 _13570_ (.A(net236),
    .B(net449),
    .X(_01703_));
 sky130_fd_sc_hd__o211a_1 _13571_ (.A1(net3221),
    .A2(net441),
    .B1(_01703_),
    .C1(net844),
    .X(_01523_));
 sky130_fd_sc_hd__or2_1 _13572_ (.A(net237),
    .B(net451),
    .X(_01704_));
 sky130_fd_sc_hd__o211a_1 _13573_ (.A1(net3325),
    .A2(net443),
    .B1(_01704_),
    .C1(net844),
    .X(_01524_));
 sky130_fd_sc_hd__or2_1 _13574_ (.A(net238),
    .B(net451),
    .X(_01705_));
 sky130_fd_sc_hd__o211a_1 _13575_ (.A1(net3323),
    .A2(net443),
    .B1(_01705_),
    .C1(net844),
    .X(_01525_));
 sky130_fd_sc_hd__or2_1 _13576_ (.A(net240),
    .B(net451),
    .X(_01706_));
 sky130_fd_sc_hd__o211a_1 _13577_ (.A1(net3462),
    .A2(net443),
    .B1(_01706_),
    .C1(net844),
    .X(_01526_));
 sky130_fd_sc_hd__or2_1 _13578_ (.A(net241),
    .B(net451),
    .X(_01707_));
 sky130_fd_sc_hd__o211a_1 _13579_ (.A1(net3455),
    .A2(net443),
    .B1(_01707_),
    .C1(net844),
    .X(_01527_));
 sky130_fd_sc_hd__nand2_1 _13580_ (.A(_01761_),
    .B(net443),
    .Y(_01708_));
 sky130_fd_sc_hd__o211a_1 _13581_ (.A1(net3466),
    .A2(net443),
    .B1(_01708_),
    .C1(net851),
    .X(_01528_));
 sky130_fd_sc_hd__or2_1 _13582_ (.A(net243),
    .B(net452),
    .X(_01709_));
 sky130_fd_sc_hd__o211a_1 _13583_ (.A1(net3468),
    .A2(net445),
    .B1(_01709_),
    .C1(net851),
    .X(_01529_));
 sky130_fd_sc_hd__or2_1 _13584_ (.A(net3394),
    .B(net452),
    .X(_01710_));
 sky130_fd_sc_hd__o211a_1 _13585_ (.A1(net3542),
    .A2(net445),
    .B1(_01710_),
    .C1(net851),
    .X(_01530_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(_01760_),
    .B(net443),
    .Y(_01711_));
 sky130_fd_sc_hd__o211a_1 _13587_ (.A1(net3522),
    .A2(net443),
    .B1(_01711_),
    .C1(net852),
    .X(_01531_));
 sky130_fd_sc_hd__or2_1 _13588_ (.A(net3368),
    .B(net451),
    .X(_01712_));
 sky130_fd_sc_hd__o211a_1 _13589_ (.A1(net3509),
    .A2(net444),
    .B1(_01712_),
    .C1(net852),
    .X(_01532_));
 sky130_fd_sc_hd__or2_1 _13590_ (.A(net3441),
    .B(net451),
    .X(_01713_));
 sky130_fd_sc_hd__o211a_1 _13591_ (.A1(net3339),
    .A2(net444),
    .B1(_01713_),
    .C1(net852),
    .X(_01533_));
 sky130_fd_sc_hd__or2_1 _13592_ (.A(net248),
    .B(net454),
    .X(_01714_));
 sky130_fd_sc_hd__o211a_1 _13593_ (.A1(net3401),
    .A2(net446),
    .B1(_01714_),
    .C1(net858),
    .X(_01534_));
 sky130_fd_sc_hd__or2_1 _13594_ (.A(net3447),
    .B(net454),
    .X(_01715_));
 sky130_fd_sc_hd__o211a_1 _13595_ (.A1(net3439),
    .A2(net446),
    .B1(_01715_),
    .C1(net858),
    .X(_01535_));
 sky130_fd_sc_hd__or2_1 _13596_ (.A(net251),
    .B(net454),
    .X(_01716_));
 sky130_fd_sc_hd__o211a_1 _13597_ (.A1(net3283),
    .A2(net446),
    .B1(_01716_),
    .C1(net858),
    .X(_01536_));
 sky130_fd_sc_hd__or2_1 _13598_ (.A(net3246),
    .B(net452),
    .X(_01717_));
 sky130_fd_sc_hd__o211a_1 _13599_ (.A1(net3184),
    .A2(net446),
    .B1(_01717_),
    .C1(net858),
    .X(_01537_));
 sky130_fd_sc_hd__o21a_1 _13600_ (.A1(net33),
    .A2(net452),
    .B1(net853),
    .X(_01538_));
 sky130_fd_sc_hd__o21a_1 _13601_ (.A1(net44),
    .A2(net452),
    .B1(net853),
    .X(_01539_));
 sky130_fd_sc_hd__or2_1 _13602_ (.A(net55),
    .B(net452),
    .X(_01718_));
 sky130_fd_sc_hd__o211a_1 _13603_ (.A1(net3211),
    .A2(net447),
    .B1(_01718_),
    .C1(net853),
    .X(_01540_));
 sky130_fd_sc_hd__and3_1 _13604_ (.A(net58),
    .B(net853),
    .C(net447),
    .X(_01541_));
 sky130_fd_sc_hd__or2_1 _13605_ (.A(net59),
    .B(net453),
    .X(_01719_));
 sky130_fd_sc_hd__o211a_1 _13606_ (.A1(net3429),
    .A2(net447),
    .B1(_01719_),
    .C1(net853),
    .X(_01542_));
 sky130_fd_sc_hd__or2_1 _13607_ (.A(net60),
    .B(net453),
    .X(_01720_));
 sky130_fd_sc_hd__o211a_1 _13608_ (.A1(net3263),
    .A2(net447),
    .B1(_01720_),
    .C1(net853),
    .X(_01543_));
 sky130_fd_sc_hd__or2_1 _13609_ (.A(net61),
    .B(net453),
    .X(_01721_));
 sky130_fd_sc_hd__o211a_1 _13610_ (.A1(net3345),
    .A2(net447),
    .B1(_01721_),
    .C1(net853),
    .X(_01544_));
 sky130_fd_sc_hd__or2_1 _13611_ (.A(net62),
    .B(net453),
    .X(_01722_));
 sky130_fd_sc_hd__o211a_1 _13612_ (.A1(net3205),
    .A2(net447),
    .B1(_01722_),
    .C1(net853),
    .X(_01545_));
 sky130_fd_sc_hd__or2_1 _13613_ (.A(net63),
    .B(net454),
    .X(_01723_));
 sky130_fd_sc_hd__o211a_1 _13614_ (.A1(net3235),
    .A2(net447),
    .B1(_01723_),
    .C1(net859),
    .X(_01546_));
 sky130_fd_sc_hd__or2_1 _13615_ (.A(net64),
    .B(net454),
    .X(_01724_));
 sky130_fd_sc_hd__o211a_1 _13616_ (.A1(net3202),
    .A2(net448),
    .B1(_01724_),
    .C1(net860),
    .X(_01547_));
 sky130_fd_sc_hd__or2_1 _13617_ (.A(net34),
    .B(net454),
    .X(_01725_));
 sky130_fd_sc_hd__o211a_1 _13618_ (.A1(net3237),
    .A2(net448),
    .B1(_01725_),
    .C1(net853),
    .X(_01548_));
 sky130_fd_sc_hd__or2_1 _13619_ (.A(net35),
    .B(net453),
    .X(_01726_));
 sky130_fd_sc_hd__o211a_1 _13620_ (.A1(net3219),
    .A2(net447),
    .B1(_01726_),
    .C1(net859),
    .X(_01549_));
 sky130_fd_sc_hd__or2_1 _13621_ (.A(net36),
    .B(net454),
    .X(_01727_));
 sky130_fd_sc_hd__o211a_1 _13622_ (.A1(net3264),
    .A2(net447),
    .B1(_01727_),
    .C1(net859),
    .X(_01550_));
 sky130_fd_sc_hd__or2_1 _13623_ (.A(net37),
    .B(net454),
    .X(_01728_));
 sky130_fd_sc_hd__o211a_1 _13624_ (.A1(net3282),
    .A2(net448),
    .B1(_01728_),
    .C1(net860),
    .X(_01551_));
 sky130_fd_sc_hd__and3_1 _13625_ (.A(net38),
    .B(net853),
    .C(net447),
    .X(_01552_));
 sky130_fd_sc_hd__or2_1 _13626_ (.A(net39),
    .B(net452),
    .X(_01729_));
 sky130_fd_sc_hd__o211a_1 _13627_ (.A1(net3464),
    .A2(net445),
    .B1(_01729_),
    .C1(net853),
    .X(_01553_));
 sky130_fd_sc_hd__or2_1 _13628_ (.A(net40),
    .B(net452),
    .X(_01730_));
 sky130_fd_sc_hd__o211a_1 _13629_ (.A1(net3226),
    .A2(net445),
    .B1(_01730_),
    .C1(net851),
    .X(_01554_));
 sky130_fd_sc_hd__or2_1 _13630_ (.A(net41),
    .B(net452),
    .X(_01731_));
 sky130_fd_sc_hd__o211a_1 _13631_ (.A1(net3496),
    .A2(net445),
    .B1(_01731_),
    .C1(net854),
    .X(_01555_));
 sky130_fd_sc_hd__or2_1 _13632_ (.A(net42),
    .B(net452),
    .X(_01732_));
 sky130_fd_sc_hd__o211a_1 _13633_ (.A1(net3536),
    .A2(net445),
    .B1(_01732_),
    .C1(net851),
    .X(_01556_));
 sky130_fd_sc_hd__or2_1 _13634_ (.A(net43),
    .B(net452),
    .X(_01733_));
 sky130_fd_sc_hd__o211a_1 _13635_ (.A1(net3495),
    .A2(net445),
    .B1(_01733_),
    .C1(net851),
    .X(_01557_));
 sky130_fd_sc_hd__or2_1 _13636_ (.A(net50),
    .B(net454),
    .X(_01734_));
 sky130_fd_sc_hd__o211a_1 _13637_ (.A1(net3392),
    .A2(net447),
    .B1(_01734_),
    .C1(net860),
    .X(_01563_));
 sky130_fd_sc_hd__or2_1 _13638_ (.A(net51),
    .B(net453),
    .X(_01735_));
 sky130_fd_sc_hd__o211a_1 _13639_ (.A1(net3452),
    .A2(net447),
    .B1(_01735_),
    .C1(net860),
    .X(_01564_));
 sky130_fd_sc_hd__or2_1 _13640_ (.A(net52),
    .B(net453),
    .X(_01736_));
 sky130_fd_sc_hd__o211a_1 _13641_ (.A1(net3420),
    .A2(net447),
    .B1(_01736_),
    .C1(net860),
    .X(_01565_));
 sky130_fd_sc_hd__or2_1 _13642_ (.A(net53),
    .B(net453),
    .X(_01737_));
 sky130_fd_sc_hd__o211a_1 _13643_ (.A1(net3421),
    .A2(net447),
    .B1(_01737_),
    .C1(net860),
    .X(_01566_));
 sky130_fd_sc_hd__or2_1 _13644_ (.A(net54),
    .B(net453),
    .X(_01738_));
 sky130_fd_sc_hd__o211a_1 _13645_ (.A1(net3461),
    .A2(net448),
    .B1(_01738_),
    .C1(net860),
    .X(_01567_));
 sky130_fd_sc_hd__or2_1 _13646_ (.A(net56),
    .B(net453),
    .X(_01739_));
 sky130_fd_sc_hd__o211a_1 _13647_ (.A1(net3435),
    .A2(net448),
    .B1(_01739_),
    .C1(net860),
    .X(_01568_));
 sky130_fd_sc_hd__or2_1 _13648_ (.A(net57),
    .B(net453),
    .X(_01740_));
 sky130_fd_sc_hd__o211a_1 _13649_ (.A1(net3216),
    .A2(net447),
    .B1(_01740_),
    .C1(net860),
    .X(_01569_));
 sky130_fd_sc_hd__nor2_4 _13650_ (.A(_02019_),
    .B(_02024_),
    .Y(_01741_));
 sky130_fd_sc_hd__mux2_1 _13651_ (.A0(net1812),
    .A1(net718),
    .S(net419),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _13652_ (.A0(net1778),
    .A1(net717),
    .S(net419),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _13653_ (.A0(net2070),
    .A1(net714),
    .S(net419),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _13654_ (.A0(net2050),
    .A1(net712),
    .S(net419),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _13655_ (.A0(net1844),
    .A1(net710),
    .S(net419),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _13656_ (.A0(net1788),
    .A1(net708),
    .S(net419),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _13657_ (.A0(net1918),
    .A1(net706),
    .S(net419),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _13658_ (.A0(net1542),
    .A1(net704),
    .S(net419),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _13659_ (.A0(net3026),
    .A1(net703),
    .S(net419),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _13660_ (.A0(net1234),
    .A1(net701),
    .S(net419),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _13661_ (.A0(net1908),
    .A1(net698),
    .S(net419),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _13662_ (.A0(net1366),
    .A1(net697),
    .S(net419),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _13663_ (.A0(net2414),
    .A1(net694),
    .S(net419),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _13664_ (.A0(net1354),
    .A1(net693),
    .S(net419),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _13665_ (.A0(net1476),
    .A1(net690),
    .S(net419),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _13666_ (.A0(net1740),
    .A1(net688),
    .S(net419),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _13667_ (.A0(net1662),
    .A1(net687),
    .S(net420),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _13668_ (.A0(net1268),
    .A1(net684),
    .S(net420),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _13669_ (.A0(net2762),
    .A1(net682),
    .S(net420),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _13670_ (.A0(net1590),
    .A1(net680),
    .S(net420),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _13671_ (.A0(net1272),
    .A1(net677),
    .S(net420),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _13672_ (.A0(net1342),
    .A1(net675),
    .S(net420),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _13673_ (.A0(net1446),
    .A1(net673),
    .S(net420),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _13674_ (.A0(net2910),
    .A1(net671),
    .S(net420),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _13675_ (.A0(net1738),
    .A1(net669),
    .S(net420),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _13676_ (.A0(net2222),
    .A1(net667),
    .S(net420),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _13677_ (.A0(net1210),
    .A1(net665),
    .S(net420),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _13678_ (.A0(net2260),
    .A1(\dpath.RF.wdata[27] ),
    .S(net420),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _13679_ (.A0(net2496),
    .A1(net661),
    .S(net420),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _13680_ (.A0(net2226),
    .A1(net658),
    .S(net420),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _13681_ (.A0(net1848),
    .A1(net657),
    .S(net420),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _13682_ (.A0(net1262),
    .A1(net655),
    .S(net420),
    .X(_01601_));
 sky130_fd_sc_hd__nor2_4 _13683_ (.A(_02019_),
    .B(_05846_),
    .Y(_01742_));
 sky130_fd_sc_hd__mux2_1 _13684_ (.A0(net2662),
    .A1(\dpath.RF.wdata[0] ),
    .S(net418),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _13685_ (.A0(net2170),
    .A1(net716),
    .S(net418),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _13686_ (.A0(net2058),
    .A1(net1374),
    .S(net418),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _13687_ (.A0(net2228),
    .A1(net713),
    .S(net418),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _13688_ (.A0(net2538),
    .A1(net711),
    .S(net418),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _13689_ (.A0(net2424),
    .A1(net709),
    .S(net418),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _13690_ (.A0(net1536),
    .A1(net707),
    .S(net418),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(net1414),
    .A1(net705),
    .S(net418),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _13692_ (.A0(net2218),
    .A1(net1180),
    .S(net418),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _13693_ (.A0(net1606),
    .A1(net701),
    .S(net418),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _13694_ (.A0(net1094),
    .A1(net1078),
    .S(net418),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _13695_ (.A0(net1672),
    .A1(net696),
    .S(net418),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _13696_ (.A0(net1698),
    .A1(net695),
    .S(net418),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _13697_ (.A0(net2738),
    .A1(net692),
    .S(net418),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _13698_ (.A0(net1804),
    .A1(net691),
    .S(net418),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _13699_ (.A0(net1504),
    .A1(net689),
    .S(net417),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _13700_ (.A0(net1300),
    .A1(net687),
    .S(net417),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _13701_ (.A0(net2116),
    .A1(net685),
    .S(net417),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _13702_ (.A0(net2502),
    .A1(net683),
    .S(net417),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _13703_ (.A0(net1774),
    .A1(net681),
    .S(net417),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _13704_ (.A0(net2614),
    .A1(net679),
    .S(net417),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _13705_ (.A0(net2708),
    .A1(net676),
    .S(net417),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _13706_ (.A0(net3052),
    .A1(net674),
    .S(net417),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _13707_ (.A0(net1574),
    .A1(net672),
    .S(net417),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _13708_ (.A0(net2364),
    .A1(net670),
    .S(net417),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _13709_ (.A0(net1314),
    .A1(net667),
    .S(net417),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _13710_ (.A0(net1714),
    .A1(net664),
    .S(net417),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _13711_ (.A0(net2554),
    .A1(net663),
    .S(net417),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _13712_ (.A0(net1702),
    .A1(net660),
    .S(net417),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _13713_ (.A0(net2660),
    .A1(net659),
    .S(net417),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _13714_ (.A0(net1678),
    .A1(net656),
    .S(net417),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _13715_ (.A0(net2150),
    .A1(net655),
    .S(_01742_),
    .X(_01633_));
 sky130_fd_sc_hd__nor2_4 _13716_ (.A(_01823_),
    .B(_01827_),
    .Y(_01743_));
 sky130_fd_sc_hd__mux2_1 _13717_ (.A0(net2556),
    .A1(net719),
    .S(net415),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _13718_ (.A0(net2392),
    .A1(net716),
    .S(net415),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _13719_ (.A0(net1530),
    .A1(net715),
    .S(net415),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _13720_ (.A0(net2564),
    .A1(net3271),
    .S(net415),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _13721_ (.A0(net1706),
    .A1(net711),
    .S(net415),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _13722_ (.A0(net1556),
    .A1(net3678),
    .S(net415),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _13723_ (.A0(net1942),
    .A1(net1360),
    .S(net415),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _13724_ (.A0(net2550),
    .A1(net704),
    .S(net415),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _13725_ (.A0(net2438),
    .A1(net702),
    .S(net415),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _13726_ (.A0(net2164),
    .A1(\dpath.RF.wdata[9] ),
    .S(net415),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _13727_ (.A0(net1660),
    .A1(net699),
    .S(net415),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _13728_ (.A0(net2928),
    .A1(net696),
    .S(net415),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _13729_ (.A0(net1850),
    .A1(net695),
    .S(net415),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _13730_ (.A0(net2028),
    .A1(net692),
    .S(net415),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _13731_ (.A0(net2290),
    .A1(net3696),
    .S(net415),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _13732_ (.A0(net1776),
    .A1(net689),
    .S(net415),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _13733_ (.A0(net1290),
    .A1(\dpath.RF.wdata[16] ),
    .S(net416),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _13734_ (.A0(net1618),
    .A1(net685),
    .S(net416),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _13735_ (.A0(net1322),
    .A1(net683),
    .S(net416),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _13736_ (.A0(net1406),
    .A1(net680),
    .S(net416),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _13737_ (.A0(net1810),
    .A1(net678),
    .S(net416),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _13738_ (.A0(net2014),
    .A1(net675),
    .S(net416),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _13739_ (.A0(net2842),
    .A1(net674),
    .S(net416),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _13740_ (.A0(net1224),
    .A1(net672),
    .S(net416),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _13741_ (.A0(net1250),
    .A1(net668),
    .S(net416),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _13742_ (.A0(net1332),
    .A1(net667),
    .S(net416),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _13743_ (.A0(net1728),
    .A1(net664),
    .S(net416),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _13744_ (.A0(net1610),
    .A1(net662),
    .S(net416),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _13745_ (.A0(net1470),
    .A1(net660),
    .S(net416),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _13746_ (.A0(net1724),
    .A1(net659),
    .S(net416),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _13747_ (.A0(net1294),
    .A1(net3712),
    .S(net416),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _13748_ (.A0(net1256),
    .A1(net654),
    .S(net416),
    .X(_01670_));
 sky130_fd_sc_hd__nor2_1 _13749_ (.A(net374),
    .B(_05991_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _13750_ (.A(net366),
    .B(_06881_),
    .Y(_01745_));
 sky130_fd_sc_hd__a2111o_1 _13751_ (.A1(net3260),
    .A2(net404),
    .B1(_02011_),
    .C1(_01744_),
    .D1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__o211a_1 _13752_ (.A1(net228),
    .A2(_02010_),
    .B1(net3261),
    .C1(net852),
    .X(_01671_));
 sky130_fd_sc_hd__o2bb2ai_1 _13753_ (.A1_N(\dpath.btarg_DX.q[1] ),
    .A2_N(net404),
    .B1(net366),
    .B2(_06882_),
    .Y(_01747_));
 sky130_fd_sc_hd__a211o_1 _13754_ (.A1(_02027_),
    .A2(_06024_),
    .B1(_01747_),
    .C1(_02011_),
    .X(_01748_));
 sky130_fd_sc_hd__o211a_1 _13755_ (.A1(net3527),
    .A2(_02010_),
    .B1(_01748_),
    .C1(net852),
    .X(_01672_));
 sky130_fd_sc_hd__clkbuf_1 _13756_ (.A(net1060),
    .X(_00769_));
 sky130_fd_sc_hd__clkbuf_1 _13757_ (.A(net1146),
    .X(_00770_));
 sky130_fd_sc_hd__clkbuf_1 _13758_ (.A(net1170),
    .X(_00771_));
 sky130_fd_sc_hd__clkbuf_1 _13759_ (.A(net1098),
    .X(_00772_));
 sky130_fd_sc_hd__clkbuf_1 _13760_ (.A(net1080),
    .X(_00773_));
 sky130_fd_sc_hd__clkbuf_1 _13761_ (.A(net1158),
    .X(_00774_));
 sky130_fd_sc_hd__clkbuf_1 _13762_ (.A(net1082),
    .X(_00775_));
 sky130_fd_sc_hd__clkbuf_1 _13763_ (.A(net1074),
    .X(_00776_));
 sky130_fd_sc_hd__clkbuf_1 _13764_ (.A(net1114),
    .X(_00777_));
 sky130_fd_sc_hd__clkbuf_1 _13765_ (.A(net1120),
    .X(_00778_));
 sky130_fd_sc_hd__clkbuf_1 _13766_ (.A(net1124),
    .X(_00779_));
 sky130_fd_sc_hd__clkbuf_1 _13767_ (.A(net1148),
    .X(_00780_));
 sky130_fd_sc_hd__clkbuf_1 _13768_ (.A(net1142),
    .X(_00781_));
 sky130_fd_sc_hd__clkbuf_1 _13769_ (.A(net1130),
    .X(_00782_));
 sky130_fd_sc_hd__clkbuf_1 _13770_ (.A(net1126),
    .X(_00783_));
 sky130_fd_sc_hd__clkbuf_1 _13771_ (.A(net1144),
    .X(_00784_));
 sky130_fd_sc_hd__clkbuf_1 _13772_ (.A(net1178),
    .X(_00785_));
 sky130_fd_sc_hd__clkbuf_1 _13773_ (.A(net1118),
    .X(_00786_));
 sky130_fd_sc_hd__clkbuf_1 _13774_ (.A(net1134),
    .X(_00787_));
 sky130_fd_sc_hd__clkbuf_1 _13775_ (.A(net1112),
    .X(_00788_));
 sky130_fd_sc_hd__clkbuf_1 _13776_ (.A(net1102),
    .X(_00789_));
 sky130_fd_sc_hd__clkbuf_1 _13777_ (.A(net1096),
    .X(_00790_));
 sky130_fd_sc_hd__clkbuf_1 _13778_ (.A(net1100),
    .X(_00791_));
 sky130_fd_sc_hd__clkbuf_1 _13779_ (.A(net1164),
    .X(_00792_));
 sky130_fd_sc_hd__clkbuf_1 _13780_ (.A(net1174),
    .X(_00793_));
 sky130_fd_sc_hd__clkbuf_1 _13781_ (.A(net1058),
    .X(_00794_));
 sky130_fd_sc_hd__clkbuf_1 _13782_ (.A(net1136),
    .X(_00795_));
 sky130_fd_sc_hd__clkbuf_1 _13783_ (.A(net1052),
    .X(_00796_));
 sky130_fd_sc_hd__clkbuf_1 _13784_ (.A(net1154),
    .X(_00797_));
 sky130_fd_sc_hd__clkbuf_1 _13785_ (.A(net1160),
    .X(_00798_));
 sky130_fd_sc_hd__clkbuf_1 _13786_ (.A(net1108),
    .X(_00799_));
 sky130_fd_sc_hd__clkbuf_1 _13787_ (.A(net1122),
    .X(_00800_));
 sky130_fd_sc_hd__o211a_1 _13788_ (.A1(net3432),
    .A2(net448),
    .B1(_05839_),
    .C1(net854),
    .X(_01558_));
 sky130_fd_sc_hd__o211a_1 _13789_ (.A1(net3393),
    .A2(net447),
    .B1(_05840_),
    .C1(net854),
    .X(_01559_));
 sky130_fd_sc_hd__o211a_1 _13790_ (.A1(net3403),
    .A2(net448),
    .B1(_05841_),
    .C1(net854),
    .X(_01560_));
 sky130_fd_sc_hd__o211a_1 _13791_ (.A1(net3285),
    .A2(net448),
    .B1(_05842_),
    .C1(net856),
    .X(_01561_));
 sky130_fd_sc_hd__o211a_1 _13792_ (.A1(net3349),
    .A2(net448),
    .B1(_05843_),
    .C1(net856),
    .X(_01562_));
 sky130_fd_sc_hd__o211a_1 _13793_ (.A1(net3464),
    .A2(net445),
    .B1(_01729_),
    .C1(net851),
    .X(_01634_));
 sky130_fd_sc_hd__o211a_1 _13794_ (.A1(net3226),
    .A2(net445),
    .B1(_01730_),
    .C1(net851),
    .X(_01635_));
 sky130_fd_sc_hd__o211a_1 _13795_ (.A1(net3496),
    .A2(net445),
    .B1(_01731_),
    .C1(net851),
    .X(_01636_));
 sky130_fd_sc_hd__o211a_1 _13796_ (.A1(net3536),
    .A2(net445),
    .B1(_01732_),
    .C1(net851),
    .X(_01637_));
 sky130_fd_sc_hd__o211a_1 _13797_ (.A1(net3495),
    .A2(net445),
    .B1(_01733_),
    .C1(net851),
    .X(_01638_));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_16_clk),
    .D(net2655),
    .Q(\dpath.RF.R[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_22_clk),
    .D(net3113),
    .Q(\dpath.RF.R[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_28_clk),
    .D(net3047),
    .Q(\dpath.RF.R[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_187_clk),
    .D(net1959),
    .Q(\dpath.RF.R[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_188_clk),
    .D(net1825),
    .Q(\dpath.RF.R[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_179_clk),
    .D(net2585),
    .Q(\dpath.RF.R[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_1_clk),
    .D(net2253),
    .Q(\dpath.RF.R[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_183_clk),
    .D(net1641),
    .Q(\dpath.RF.R[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_28_clk),
    .D(net2831),
    .Q(\dpath.RF.R[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_156_clk),
    .D(net2103),
    .Q(\dpath.RF.R[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_149_clk),
    .D(net2433),
    .Q(\dpath.RF.R[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_176_clk),
    .D(net2967),
    .Q(\dpath.RF.R[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_159_clk),
    .D(net2201),
    .Q(\dpath.RF.R[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_173_clk),
    .D(net2211),
    .Q(\dpath.RF.R[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_161_clk),
    .D(net2225),
    .Q(\dpath.RF.R[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_166_clk),
    .D(net2447),
    .Q(\dpath.RF.R[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_123_clk),
    .D(net1931),
    .Q(\dpath.RF.R[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_167_clk),
    .D(net2157),
    .Q(\dpath.RF.R[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_117_clk),
    .D(net2697),
    .Q(\dpath.RF.R[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_163_clk),
    .D(net2133),
    .Q(\dpath.RF.R[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_116_clk),
    .D(net2927),
    .Q(\dpath.RF.R[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_108_clk),
    .D(net2391),
    .Q(\dpath.RF.R[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_151_clk),
    .D(net2657),
    .Q(\dpath.RF.R[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_128_clk),
    .D(net1763),
    .Q(\dpath.RF.R[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_111_clk),
    .D(net2377),
    .Q(\dpath.RF.R[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_83_clk),
    .D(net1657),
    .Q(\dpath.RF.R[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_150_clk),
    .D(net3089),
    .Q(\dpath.RF.R[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_84_clk),
    .D(net3131),
    .Q(\dpath.RF.R[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_136_clk),
    .D(net2849),
    .Q(\dpath.RF.R[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_77_clk),
    .D(net1897),
    .Q(\dpath.RF.R[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_141_clk),
    .D(net1915),
    .Q(\dpath.RF.R[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_77_clk),
    .D(net2305),
    .Q(\dpath.RF.R[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_16_clk),
    .D(net2865),
    .Q(\dpath.RF.R[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_22_clk),
    .D(net1651),
    .Q(\dpath.RF.R[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_34_clk),
    .D(net1755),
    .Q(\dpath.RF.R[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_187_clk),
    .D(net2321),
    .Q(\dpath.RF.R[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_188_clk),
    .D(net1705),
    .Q(\dpath.RF.R[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_179_clk),
    .D(net1921),
    .Q(\dpath.RF.R[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_188_clk),
    .D(net1925),
    .Q(\dpath.RF.R[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_186_clk),
    .D(net3041),
    .Q(\dpath.RF.R[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_28_clk),
    .D(net1801),
    .Q(\dpath.RF.R[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_156_clk),
    .D(net2597),
    .Q(\dpath.RF.R[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_149_clk),
    .D(net1985),
    .Q(\dpath.RF.R[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_176_clk),
    .D(net1583),
    .Q(\dpath.RF.R[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_159_clk),
    .D(net2775),
    .Q(\dpath.RF.R[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_173_clk),
    .D(net2917),
    .Q(\dpath.RF.R[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_161_clk),
    .D(net2465),
    .Q(\dpath.RF.R[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_172_clk),
    .D(net2665),
    .Q(\dpath.RF.R[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_123_clk),
    .D(net2197),
    .Q(\dpath.RF.R[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_167_clk),
    .D(net2895),
    .Q(\dpath.RF.R[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_117_clk),
    .D(net1559),
    .Q(\dpath.RF.R[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_163_clk),
    .D(net1461),
    .Q(\dpath.RF.R[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_116_clk),
    .D(net1555),
    .Q(\dpath.RF.R[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_115_clk),
    .D(net1293),
    .Q(\dpath.RF.R[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_151_clk),
    .D(net2173),
    .Q(\dpath.RF.R[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_128_clk),
    .D(net1581),
    .Q(\dpath.RF.R[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_111_clk),
    .D(net2235),
    .Q(\dpath.RF.R[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_133_clk),
    .D(net1635),
    .Q(\dpath.RF.R[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_150_clk),
    .D(net2553),
    .Q(\dpath.RF.R[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_81_clk),
    .D(net2583),
    .Q(\dpath.RF.R[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_136_clk),
    .D(net2035),
    .Q(\dpath.RF.R[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_77_clk),
    .D(net1841),
    .Q(\dpath.RF.R[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_141_clk),
    .D(net2941),
    .Q(\dpath.RF.R[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_77_clk),
    .D(net1767),
    .Q(\dpath.RF.R[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_16_clk),
    .D(net2999),
    .Q(\dpath.RF.R[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_23_clk),
    .D(net2549),
    .Q(\dpath.RF.R[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_28_clk),
    .D(net2945),
    .Q(\dpath.RF.R[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_181_clk),
    .D(net3071),
    .Q(\dpath.RF.R[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_1_clk),
    .D(net2647),
    .Q(\dpath.RF.R[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_179_clk),
    .D(net2385),
    .Q(\dpath.RF.R[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_1_clk),
    .D(net2893),
    .Q(\dpath.RF.R[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_184_clk),
    .D(net2785),
    .Q(\dpath.RF.R[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_34_clk),
    .D(net2003),
    .Q(\dpath.RF.R[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_155_clk),
    .D(net2735),
    .Q(\dpath.RF.R[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_149_clk),
    .D(net2317),
    .Q(\dpath.RF.R[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_176_clk),
    .D(net2719),
    .Q(\dpath.RF.R[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_159_clk),
    .D(net3075),
    .Q(\dpath.RF.R[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_173_clk),
    .D(net2095),
    .Q(\dpath.RF.R[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_161_clk),
    .D(net2755),
    .Q(\dpath.RF.R[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_166_clk),
    .D(net2641),
    .Q(\dpath.RF.R[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_123_clk),
    .D(net2685),
    .Q(\dpath.RF.R[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_122_clk),
    .D(net2619),
    .Q(\dpath.RF.R[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_117_clk),
    .D(net2987),
    .Q(\dpath.RF.R[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_126_clk),
    .D(net2183),
    .Q(\dpath.RF.R[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_115_clk),
    .D(net2283),
    .Q(\dpath.RF.R[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_109_clk),
    .D(net2277),
    .Q(\dpath.RF.R[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_139_clk),
    .D(net1941),
    .Q(\dpath.RF.R[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_131_clk),
    .D(net3049),
    .Q(\dpath.RF.R[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_111_clk),
    .D(net2789),
    .Q(\dpath.RF.R[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_103_clk),
    .D(net3151),
    .Q(\dpath.RF.R[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_150_clk),
    .D(net3193),
    .Q(\dpath.RF.R[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_84_clk),
    .D(net2233),
    .Q(\dpath.RF.R[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_79_clk),
    .D(net2245),
    .Q(\dpath.RF.R[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_87_clk),
    .D(net2809),
    .Q(\dpath.RF.R[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_142_clk),
    .D(net2765),
    .Q(\dpath.RF.R[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_87_clk),
    .D(net2713),
    .Q(\dpath.RF.R[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_23_clk),
    .D(net2745),
    .Q(\dpath.RF.R[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_24_clk),
    .D(net2487),
    .Q(\dpath.RF.R[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_30_clk),
    .D(net3011),
    .Q(\dpath.RF.R[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_180_clk),
    .D(net3083),
    .Q(\dpath.RF.R[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_2_clk),
    .D(net2459),
    .Q(\dpath.RF.R[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_158_clk),
    .D(net3105),
    .Q(\dpath.RF.R[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_2_clk),
    .D(net3043),
    .Q(\dpath.RF.R[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_180_clk),
    .D(net2953),
    .Q(\dpath.RF.R[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_33_clk),
    .D(net3183),
    .Q(\dpath.RF.R[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_154_clk),
    .D(net2959),
    .Q(\dpath.RF.R[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_148_clk),
    .D(net2625),
    .Q(\dpath.RF.R[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_177_clk),
    .D(net3169),
    .Q(\dpath.RF.R[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_163_clk),
    .D(net2991),
    .Q(\dpath.RF.R[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_160_clk),
    .D(net2955),
    .Q(\dpath.RF.R[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_152_clk),
    .D(net2977),
    .Q(\dpath.RF.R[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_164_clk),
    .D(net2577),
    .Q(\dpath.RF.R[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_124_clk),
    .D(net2445),
    .Q(\dpath.RF.R[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_126_clk),
    .D(net2689),
    .Q(\dpath.RF.R[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_130_clk),
    .D(net2563),
    .Q(\dpath.RF.R[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_127_clk),
    .D(net2837),
    .Q(\dpath.RF.R[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_113_clk),
    .D(net2771),
    .Q(\dpath.RF.R[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_112_clk),
    .D(net2595),
    .Q(\dpath.RF.R[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_138_clk),
    .D(net3081),
    .Q(\dpath.RF.R[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_135_clk),
    .D(net2639),
    .Q(\dpath.RF.R[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_132_clk),
    .D(net3013),
    .Q(\dpath.RF.R[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_133_clk),
    .D(net3175),
    .Q(\dpath.RF.R[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_145_clk),
    .D(net3107),
    .Q(\dpath.RF.R[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_81_clk),
    .D(net3145),
    .Q(\dpath.RF.R[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_73_clk),
    .D(net3031),
    .Q(\dpath.RF.R[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_76_clk),
    .D(net2703),
    .Q(\dpath.RF.R[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_143_clk),
    .D(net3077),
    .Q(\dpath.RF.R[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_77_clk),
    .D(net2899),
    .Q(\dpath.RF.R[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_23_clk),
    .D(net3181),
    .Q(\dpath.RF.R[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_24_clk),
    .D(net2613),
    .Q(\dpath.RF.R[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_32_clk),
    .D(net1871),
    .Q(\dpath.RF.R[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_180_clk),
    .D(net2901),
    .Q(\dpath.RF.R[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_179_clk),
    .D(net2629),
    .Q(\dpath.RF.R[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_158_clk),
    .D(net2701),
    .Q(\dpath.RF.R[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_179_clk),
    .D(net2607),
    .Q(\dpath.RF.R[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_178_clk),
    .D(net3029),
    .Q(\dpath.RF.R[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_36_clk),
    .D(net2921),
    .Q(\dpath.RF.R[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_154_clk),
    .D(net2875),
    .Q(\dpath.RF.R[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_147_clk),
    .D(net2971),
    .Q(\dpath.RF.R[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_177_clk),
    .D(net3173),
    .Q(\dpath.RF.R[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_162_clk),
    .D(net3103),
    .Q(\dpath.RF.R[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_160_clk),
    .D(net3141),
    .Q(\dpath.RF.R[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_151_clk),
    .D(net3127),
    .Q(\dpath.RF.R[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_163_clk),
    .D(net2915),
    .Q(\dpath.RF.R[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_129_clk),
    .D(net3079),
    .Q(\dpath.RF.R[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_125_clk),
    .D(net3021),
    .Q(\dpath.RF.R[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_131_clk),
    .D(net3125),
    .Q(\dpath.RF.R[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_129_clk),
    .D(net2979),
    .Q(\dpath.RF.R[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_112_clk),
    .D(net2711),
    .Q(\dpath.RF.R[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_112_clk),
    .D(net2985),
    .Q(\dpath.RF.R[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_137_clk),
    .D(net2195),
    .Q(\dpath.RF.R[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_134_clk),
    .D(net2861),
    .Q(\dpath.RF.R[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_133_clk),
    .D(net2573),
    .Q(\dpath.RF.R[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_82_clk),
    .D(net2617),
    .Q(\dpath.RF.R[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13952_ (.CLK(clknet_leaf_145_clk),
    .D(net2467),
    .Q(\dpath.RF.R[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13953_ (.CLK(clknet_leaf_81_clk),
    .D(net3129),
    .Q(\dpath.RF.R[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_74_clk),
    .D(net2853),
    .Q(\dpath.RF.R[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13955_ (.CLK(clknet_leaf_76_clk),
    .D(net2637),
    .Q(\dpath.RF.R[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13956_ (.CLK(clknet_leaf_72_clk),
    .D(net2375),
    .Q(\dpath.RF.R[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13957_ (.CLK(clknet_leaf_77_clk),
    .D(net2239),
    .Q(\dpath.RF.R[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13958_ (.CLK(clknet_leaf_21_clk),
    .D(net3153),
    .Q(\dpath.RF.R[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13959_ (.CLK(clknet_leaf_4_clk),
    .D(net2839),
    .Q(\dpath.RF.R[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13960_ (.CLK(clknet_leaf_30_clk),
    .D(net2443),
    .Q(\dpath.RF.R[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13961_ (.CLK(clknet_leaf_187_clk),
    .D(net2421),
    .Q(\dpath.RF.R[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13962_ (.CLK(clknet_leaf_188_clk),
    .D(net2815),
    .Q(\dpath.RF.R[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13963_ (.CLK(clknet_leaf_178_clk),
    .D(net3119),
    .Q(\dpath.RF.R[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13964_ (.CLK(clknet_leaf_188_clk),
    .D(net3187),
    .Q(\dpath.RF.R[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13965_ (.CLK(clknet_leaf_186_clk),
    .D(net2355),
    .Q(\dpath.RF.R[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13966_ (.CLK(clknet_leaf_34_clk),
    .D(net2645),
    .Q(\dpath.RF.R[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13967_ (.CLK(clknet_leaf_156_clk),
    .D(net2797),
    .Q(\dpath.RF.R[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13968_ (.CLK(clknet_leaf_35_clk),
    .D(net2419),
    .Q(\dpath.RF.R[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13969_ (.CLK(clknet_leaf_175_clk),
    .D(net2795),
    .Q(\dpath.RF.R[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13970_ (.CLK(clknet_leaf_158_clk),
    .D(net2257),
    .Q(\dpath.RF.R[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13971_ (.CLK(clknet_leaf_172_clk),
    .D(net2509),
    .Q(\dpath.RF.R[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13972_ (.CLK(clknet_leaf_153_clk),
    .D(net1969),
    .Q(\dpath.RF.R[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13973_ (.CLK(clknet_leaf_171_clk),
    .D(net2215),
    .Q(\dpath.RF.R[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13974_ (.CLK(clknet_leaf_122_clk),
    .D(net2975),
    .Q(\dpath.RF.R[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13975_ (.CLK(clknet_leaf_168_clk),
    .D(net2523),
    .Q(\dpath.RF.R[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13976_ (.CLK(clknet_leaf_118_clk),
    .D(net2743),
    .Q(\dpath.RF.R[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13977_ (.CLK(clknet_leaf_162_clk),
    .D(net2897),
    .Q(\dpath.RF.R[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_116_clk),
    .D(net3121),
    .Q(\dpath.RF.R[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_109_clk),
    .D(net2671),
    .Q(\dpath.RF.R[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_140_clk),
    .D(net2559),
    .Q(\dpath.RF.R[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_128_clk),
    .D(net2751),
    .Q(\dpath.RF.R[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_110_clk),
    .D(net2535),
    .Q(\dpath.RF.R[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_103_clk),
    .D(net2769),
    .Q(\dpath.RF.R[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_148_clk),
    .D(net2675),
    .Q(\dpath.RF.R[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_84_clk),
    .D(net2073),
    .Q(\dpath.RF.R[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_79_clk),
    .D(net2299),
    .Q(\dpath.RF.R[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_78_clk),
    .D(net2827),
    .Q(\dpath.RF.R[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_141_clk),
    .D(net2403),
    .Q(\dpath.RF.R[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_88_clk),
    .D(net2511),
    .Q(\dpath.RF.R[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_16_clk),
    .D(net2933),
    .Q(\dpath.RF.R[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_23_clk),
    .D(net2543),
    .Q(\dpath.RF.R[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_29_clk),
    .D(net1997),
    .Q(\dpath.RF.R[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_182_clk),
    .D(net1577),
    .Q(\dpath.RF.R[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_1_clk),
    .D(net2049),
    .Q(\dpath.RF.R[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_179_clk),
    .D(net1283),
    .Q(\dpath.RF.R[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_1_clk),
    .D(net2783),
    .Q(\dpath.RF.R[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_185_clk),
    .D(net1613),
    .Q(\dpath.RF.R[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_28_clk),
    .D(net1317),
    .Q(\dpath.RF.R[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_155_clk),
    .D(net2601),
    .Q(\dpath.RF.R[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_149_clk),
    .D(net2721),
    .Q(\dpath.RF.R[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_176_clk),
    .D(net1787),
    .Q(\dpath.RF.R[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_159_clk),
    .D(net1199),
    .Q(\dpath.RF.R[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14003_ (.CLK(clknet_leaf_173_clk),
    .D(net2867),
    .Q(\dpath.RF.R[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_161_clk),
    .D(net2749),
    .Q(\dpath.RF.R[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_166_clk),
    .D(net1609),
    .Q(\dpath.RF.R[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_123_clk),
    .D(net2339),
    .Q(\dpath.RF.R[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_167_clk),
    .D(net1187),
    .Q(\dpath.RF.R[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_117_clk),
    .D(net1951),
    .Q(\dpath.RF.R[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_126_clk),
    .D(net2331),
    .Q(\dpath.RF.R[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_115_clk),
    .D(net1513),
    .Q(\dpath.RF.R[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_109_clk),
    .D(net1517),
    .Q(\dpath.RF.R[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_151_clk),
    .D(net1571),
    .Q(\dpath.RF.R[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_131_clk),
    .D(net1735),
    .Q(\dpath.RF.R[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_111_clk),
    .D(net2031),
    .Q(\dpath.RF.R[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_103_clk),
    .D(net2399),
    .Q(\dpath.RF.R[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_150_clk),
    .D(net3167),
    .Q(\dpath.RF.R[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_84_clk),
    .D(net1671),
    .Q(\dpath.RF.R[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_79_clk),
    .D(net1189),
    .Q(\dpath.RF.R[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_87_clk),
    .D(net2347),
    .Q(\dpath.RF.R[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_141_clk),
    .D(net1297),
    .Q(\dpath.RF.R[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_87_clk),
    .D(net2043),
    .Q(\dpath.RF.R[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_13_clk),
    .D(_00234_),
    .Q(\ctrl.val_D ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_43_clk),
    .D(net3199),
    .Q(\ctrl.val_MW.q ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_48_clk),
    .D(net1177),
    .Q(\ctrl.inst_M[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_53_clk),
    .D(net1209),
    .Q(\ctrl.inst_M[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_48_clk),
    .D(net1167),
    .Q(\ctrl.inst_M[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_47_clk),
    .D(net1151),
    .Q(\ctrl.inst_M[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_47_clk),
    .D(_00240_),
    .Q(\ctrl.inst_M[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_47_clk),
    .D(_00241_),
    .Q(\ctrl.inst_M[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_47_clk),
    .D(net1469),
    .Q(\ctrl.inst_M[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_45_clk),
    .D(_00243_),
    .Q(\ctrl.inst_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_43_clk),
    .D(_00244_),
    .Q(\ctrl.inst_M[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_45_clk),
    .D(_00245_),
    .Q(\ctrl.inst_M[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_46_clk),
    .D(_00246_),
    .Q(\ctrl.inst_M[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_46_clk),
    .D(_00247_),
    .Q(\ctrl.inst_M[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_47_clk),
    .D(_00248_),
    .Q(\ctrl.inst_M[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_47_clk),
    .D(net2869),
    .Q(\ctrl.inst_M[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_47_clk),
    .D(net2973),
    .Q(\ctrl.inst_M[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_66_clk),
    .D(_00251_),
    .Q(\ctrl.inst_M[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_67_clk),
    .D(_00252_),
    .Q(\ctrl.inst_M[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_67_clk),
    .D(_00253_),
    .Q(\ctrl.inst_M[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_67_clk),
    .D(_00254_),
    .Q(\ctrl.inst_M[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_43_clk),
    .D(net1001),
    .Q(\ctrl.inst_M[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_42_clk),
    .D(net1093),
    .Q(\ctrl.inst_M[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_42_clk),
    .D(net991),
    .Q(\ctrl.inst_M[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_42_clk),
    .D(net911),
    .Q(\ctrl.inst_M[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_42_clk),
    .D(net907),
    .Q(\ctrl.inst_M[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_42_clk),
    .D(net915),
    .Q(\ctrl.inst_M[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_42_clk),
    .D(net913),
    .Q(\ctrl.inst_M[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_47_clk),
    .D(net1091),
    .Q(\ctrl.inst_M[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_49_clk),
    .D(_00263_),
    .Q(\ctrl.val_DX.q ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_50_clk),
    .D(net2061),
    .Q(\ctrl.inst_X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_50_clk),
    .D(net2407),
    .Q(\ctrl.inst_X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_51_clk),
    .D(_00266_),
    .Q(\ctrl.inst_X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_51_clk),
    .D(net3177),
    .Q(\ctrl.inst_X[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_53_clk),
    .D(_00268_),
    .Q(\ctrl.inst_X[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_53_clk),
    .D(_00269_),
    .Q(\ctrl.inst_X[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_53_clk),
    .D(_00270_),
    .Q(\ctrl.inst_X[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_48_clk),
    .D(_00271_),
    .Q(\ctrl.inst_X[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_48_clk),
    .D(_00272_),
    .Q(\ctrl.inst_X[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_48_clk),
    .D(_00273_),
    .Q(\ctrl.inst_X[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_46_clk),
    .D(_00274_),
    .Q(\ctrl.inst_X[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_46_clk),
    .D(_00275_),
    .Q(\ctrl.inst_X[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_53_clk),
    .D(_00276_),
    .Q(\ctrl.inst_X[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_53_clk),
    .D(_00277_),
    .Q(\ctrl.inst_X[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_53_clk),
    .D(_00278_),
    .Q(\ctrl.inst_X[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_40_clk),
    .D(_00279_),
    .Q(\ctrl.inst_X[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_41_clk),
    .D(_00280_),
    .Q(\ctrl.inst_X[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_40_clk),
    .D(_00281_),
    .Q(\ctrl.inst_X[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_41_clk),
    .D(_00282_),
    .Q(\ctrl.inst_X[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_43_clk),
    .D(_00283_),
    .Q(\ctrl.inst_X[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_53_clk),
    .D(_00284_),
    .Q(\ctrl.inst_X[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_54_clk),
    .D(_00285_),
    .Q(\ctrl.inst_X[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_56_clk),
    .D(_00286_),
    .Q(\ctrl.inst_X[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_56_clk),
    .D(_00287_),
    .Q(\ctrl.inst_X[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_54_clk),
    .D(_00288_),
    .Q(\ctrl.inst_X[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_56_clk),
    .D(_00289_),
    .Q(\ctrl.inst_X[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_54_clk),
    .D(_00290_),
    .Q(\ctrl.inst_X[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_47_clk),
    .D(net1023),
    .Q(\ctrl.inst_W[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_48_clk),
    .D(net973),
    .Q(\ctrl.inst_W[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_43_clk),
    .D(_00293_),
    .Q(\ctrl.inst_W[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14082_ (.CLK(clknet_leaf_46_clk),
    .D(net3213),
    .Q(\ctrl.inst_W[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_47_clk),
    .D(_00295_),
    .Q(\ctrl.inst_W[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_42_clk),
    .D(_00296_),
    .Q(\ctrl.inst_W[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_42_clk),
    .D(net3117),
    .Q(\ctrl.inst_W[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14086_ (.CLK(clknet_leaf_44_clk),
    .D(_00298_),
    .Q(\ctrl.c2d_rf_waddr_W[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14087_ (.CLK(clknet_leaf_44_clk),
    .D(_00299_),
    .Q(\ctrl.c2d_rf_waddr_W[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14088_ (.CLK(clknet_leaf_43_clk),
    .D(_00300_),
    .Q(\ctrl.c2d_rf_waddr_W[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14089_ (.CLK(clknet_leaf_44_clk),
    .D(_00301_),
    .Q(\ctrl.c2d_rf_waddr_W[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14090_ (.CLK(clknet_leaf_43_clk),
    .D(_00302_),
    .Q(\ctrl.c2d_rf_waddr_W[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_42_clk),
    .D(net3087),
    .Q(\ctrl.inst_W[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_42_clk),
    .D(net1133),
    .Q(\ctrl.inst_W[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_42_clk),
    .D(net1169),
    .Q(\ctrl.inst_W[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14094_ (.CLK(clknet_leaf_65_clk),
    .D(net945),
    .Q(\ctrl.inst_W[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_66_clk),
    .D(net925),
    .Q(\ctrl.inst_W[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_66_clk),
    .D(net933),
    .Q(\ctrl.inst_W[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_66_clk),
    .D(net923),
    .Q(\ctrl.inst_W[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_43_clk),
    .D(net1007),
    .Q(\ctrl.inst_W[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_42_clk),
    .D(net1041),
    .Q(\ctrl.inst_W[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_42_clk),
    .D(net1217),
    .Q(\ctrl.inst_W[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_42_clk),
    .D(net1153),
    .Q(\ctrl.inst_W[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_42_clk),
    .D(net1117),
    .Q(\ctrl.inst_W[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_42_clk),
    .D(net1139),
    .Q(\ctrl.inst_W[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_42_clk),
    .D(net1163),
    .Q(\ctrl.inst_W[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_42_clk),
    .D(net961),
    .Q(\ctrl.inst_W[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_20_clk),
    .D(net1881),
    .Q(\dpath.RF.R[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_26_clk),
    .D(net1791),
    .Q(\dpath.RF.R[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_31_clk),
    .D(net1413),
    .Q(\dpath.RF.R[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_183_clk),
    .D(net1923),
    .Q(\dpath.RF.R[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_180_clk),
    .D(net2323),
    .Q(\dpath.RF.R[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_156_clk),
    .D(net2009),
    .Q(\dpath.RF.R[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_24_clk),
    .D(net2427),
    .Q(\dpath.RF.R[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14113_ (.CLK(clknet_leaf_184_clk),
    .D(net1989),
    .Q(\dpath.RF.R[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_33_clk),
    .D(net1181),
    .Q(\dpath.RF.R[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_154_clk),
    .D(net2349),
    .Q(\dpath.RF.R[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14116_ (.CLK(clknet_leaf_37_clk),
    .D(net1457),
    .Q(\dpath.RF.R[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_177_clk),
    .D(net2747),
    .Q(\dpath.RF.R[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_161_clk),
    .D(net2423),
    .Q(\dpath.RF.R[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14119_ (.CLK(clknet_leaf_172_clk),
    .D(net2623),
    .Q(\dpath.RF.R[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14120_ (.CLK(clknet_leaf_151_clk),
    .D(net2707),
    .Q(\dpath.RF.R[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_166_clk),
    .D(net1753),
    .Q(\dpath.RF.R[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_123_clk),
    .D(net1979),
    .Q(\dpath.RF.R[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_122_clk),
    .D(net2589),
    .Q(\dpath.RF.R[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_118_clk),
    .D(net2065),
    .Q(\dpath.RF.R[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_128_clk),
    .D(net2643),
    .Q(\dpath.RF.R[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_115_clk),
    .D(net1837),
    .Q(\dpath.RF.R[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_112_clk),
    .D(net2759),
    .Q(\dpath.RF.R[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_137_clk),
    .D(net2567),
    .Q(\dpath.RF.R[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_136_clk),
    .D(net2939),
    .Q(\dpath.RF.R[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_111_clk),
    .D(net2579),
    .Q(\dpath.RF.R[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_82_clk),
    .D(net2371),
    .Q(\dpath.RF.R[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_147_clk),
    .D(net1903),
    .Q(\dpath.RF.R[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_80_clk),
    .D(net1655),
    .Q(\dpath.RF.R[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_69_clk),
    .D(net2521),
    .Q(\dpath.RF.R[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_68_clk),
    .D(net2135),
    .Q(\dpath.RF.R[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_71_clk),
    .D(net2803),
    .Q(\dpath.RF.R[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_76_clk),
    .D(net2817),
    .Q(\dpath.RF.R[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_20_clk),
    .D(net1287),
    .Q(\dpath.RF.R[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_26_clk),
    .D(net1899),
    .Q(\dpath.RF.R[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_31_clk),
    .D(net3001),
    .Q(\dpath.RF.R[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_182_clk),
    .D(net1255),
    .Q(\dpath.RF.R[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_181_clk),
    .D(net1647),
    .Q(\dpath.RF.R[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_179_clk),
    .D(net2575),
    .Q(\dpath.RF.R[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_3_clk),
    .D(net3189),
    .Q(\dpath.RF.R[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_184_clk),
    .D(net2129),
    .Q(\dpath.RF.R[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_39_clk),
    .D(net2723),
    .Q(\dpath.RF.R[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_26_clk),
    .D(net2825),
    .Q(\dpath.RF.R[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_36_clk),
    .D(net1795),
    .Q(\dpath.RF.R[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_176_clk),
    .D(net2541),
    .Q(\dpath.RF.R[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_161_clk),
    .D(net1451),
    .Q(\dpath.RF.R[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_177_clk),
    .D(net1961),
    .Q(\dpath.RF.R[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_154_clk),
    .D(net1597),
    .Q(\dpath.RF.R[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_165_clk),
    .D(net1501),
    .Q(\dpath.RF.R[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_123_clk),
    .D(net2011),
    .Q(\dpath.RF.R[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_164_clk),
    .D(net1065),
    .Q(\dpath.RF.R[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_130_clk),
    .D(net1201),
    .Q(\dpath.RF.R[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_127_clk),
    .D(net1313),
    .Q(\dpath.RF.R[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_114_clk),
    .D(net1411),
    .Q(\dpath.RF.R[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_113_clk),
    .D(net1285),
    .Q(\dpath.RF.R[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_139_clk),
    .D(net1587),
    .Q(\dpath.RF.R[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_137_clk),
    .D(net1541),
    .Q(\dpath.RF.R[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_132_clk),
    .D(net1363),
    .Q(\dpath.RF.R[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_133_clk),
    .D(net1373),
    .Q(\dpath.RF.R[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_147_clk),
    .D(net2495),
    .Q(\dpath.RF.R[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_79_clk),
    .D(net1529),
    .Q(\dpath.RF.R[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_69_clk),
    .D(net1389),
    .Q(\dpath.RF.R[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_69_clk),
    .D(net1721),
    .Q(\dpath.RF.R[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_145_clk),
    .D(net1253),
    .Q(\dpath.RF.R[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_75_clk),
    .D(net2131),
    .Q(\dpath.RF.R[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_175_clk),
    .D(net1069),
    .Q(net196));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_174_clk),
    .D(net909),
    .Q(net207));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_174_clk),
    .D(net1085),
    .Q(net218));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_175_clk),
    .D(net1107),
    .Q(net221));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_175_clk),
    .D(net1129),
    .Q(net222));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_174_clk),
    .D(net1111),
    .Q(net223));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_170_clk),
    .D(net1071),
    .Q(net224));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_170_clk),
    .D(net987),
    .Q(net225));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_170_clk),
    .D(net1047),
    .Q(net226));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_174_clk),
    .D(net1027),
    .Q(net227));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_170_clk),
    .D(_00392_),
    .Q(net197));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_169_clk),
    .D(net1031),
    .Q(net198));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_169_clk),
    .D(net1025),
    .Q(net199));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_169_clk),
    .D(net1045),
    .Q(net200));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_169_clk),
    .D(net1039),
    .Q(net201));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_169_clk),
    .D(net1021),
    .Q(net202));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_121_clk),
    .D(net1073),
    .Q(net203));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_121_clk),
    .D(net1015),
    .Q(net204));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_120_clk),
    .D(net1087),
    .Q(net205));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_120_clk),
    .D(net1035),
    .Q(net206));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_120_clk),
    .D(net1077),
    .Q(net208));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_120_clk),
    .D(net1105),
    .Q(net209));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_120_clk),
    .D(net1089),
    .Q(net210));
 sky130_fd_sc_hd__dfxtp_1 _14193_ (.CLK(clknet_leaf_119_clk),
    .D(net1051),
    .Q(net211));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_119_clk),
    .D(net1057),
    .Q(net212));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_119_clk),
    .D(net1063),
    .Q(net213));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_120_clk),
    .D(_00408_),
    .Q(net214));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_119_clk),
    .D(_00409_),
    .Q(net215));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_117_clk),
    .D(_00410_),
    .Q(net216));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_117_clk),
    .D(_00411_),
    .Q(net217));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_117_clk),
    .D(_00412_),
    .Q(net219));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_117_clk),
    .D(_00413_),
    .Q(net220));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_20_clk),
    .D(net2079),
    .Q(\dpath.RF.R[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_25_clk),
    .D(net1393),
    .Q(\dpath.RF.R[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_31_clk),
    .D(net2533),
    .Q(\dpath.RF.R[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_183_clk),
    .D(net2635),
    .Q(\dpath.RF.R[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_180_clk),
    .D(net2381),
    .Q(\dpath.RF.R[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_179_clk),
    .D(net2591),
    .Q(\dpath.RF.R[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_3_clk),
    .D(net2989),
    .Q(\dpath.RF.R[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_184_clk),
    .D(net1697),
    .Q(\dpath.RF.R[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_32_clk),
    .D(net1391),
    .Q(\dpath.RF.R[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_27_clk),
    .D(net1473),
    .Q(\dpath.RF.R[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_36_clk),
    .D(net1945),
    .Q(\dpath.RF.R[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_176_clk),
    .D(net2561),
    .Q(\dpath.RF.R[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_161_clk),
    .D(net2829),
    .Q(\dpath.RF.R[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_172_clk),
    .D(net2039),
    .Q(\dpath.RF.R[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_149_clk),
    .D(net2965),
    .Q(\dpath.RF.R[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_165_clk),
    .D(net2363),
    .Q(\dpath.RF.R[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14218_ (.CLK(clknet_leaf_125_clk),
    .D(net1907),
    .Q(\dpath.RF.R[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_167_clk),
    .D(net2099),
    .Q(\dpath.RF.R[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_130_clk),
    .D(net2801),
    .Q(\dpath.RF.R[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_138_clk),
    .D(net999),
    .Q(\dpath.RF.R[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_114_clk),
    .D(net2319),
    .Q(\dpath.RF.R[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_112_clk),
    .D(net2599),
    .Q(\dpath.RF.R[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_138_clk),
    .D(net3061),
    .Q(\dpath.RF.R[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_137_clk),
    .D(net2189),
    .Q(\dpath.RF.R[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_112_clk),
    .D(net3101),
    .Q(\dpath.RF.R[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_133_clk),
    .D(net2353),
    .Q(\dpath.RF.R[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_147_clk),
    .D(net2517),
    .Q(\dpath.RF.R[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_80_clk),
    .D(net2493),
    .Q(\dpath.RF.R[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_75_clk),
    .D(net1731),
    .Q(\dpath.RF.R[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_76_clk),
    .D(net3009),
    .Q(\dpath.RF.R[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_146_clk),
    .D(net1719),
    .Q(\dpath.RF.R[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_76_clk),
    .D(net2361),
    .Q(\dpath.RF.R[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_23_clk),
    .D(net2925),
    .Q(\dpath.RF.R[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_26_clk),
    .D(net2981),
    .Q(\dpath.RF.R[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_31_clk),
    .D(net1223),
    .Q(\dpath.RF.R[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_180_clk),
    .D(net2727),
    .Q(\dpath.RF.R[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_180_clk),
    .D(net2413),
    .Q(\dpath.RF.R[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_156_clk),
    .D(net2887),
    .Q(\dpath.RF.R[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_24_clk),
    .D(net1809),
    .Q(\dpath.RF.R[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_176_clk),
    .D(net2263),
    .Q(\dpath.RF.R[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_37_clk),
    .D(net1629),
    .Q(\dpath.RF.R[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_154_clk),
    .D(net2287),
    .Q(\dpath.RF.R[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_38_clk),
    .D(net1727),
    .Q(\dpath.RF.R[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_177_clk),
    .D(net1869),
    .Q(\dpath.RF.R[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_162_clk),
    .D(net2715),
    .Q(\dpath.RF.R[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_165_clk),
    .D(net2731),
    .Q(\dpath.RF.R[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_151_clk),
    .D(net2821),
    .Q(\dpath.RF.R[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_164_clk),
    .D(net1497),
    .Q(\dpath.RF.R[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_118_clk),
    .D(net1441),
    .Q(\dpath.RF.R[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_122_clk),
    .D(net1957),
    .Q(\dpath.RF.R[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_114_clk),
    .D(net2603),
    .Q(\dpath.RF.R[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_138_clk),
    .D(net2329),
    .Q(\dpath.RF.R[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_115_clk),
    .D(net1429),
    .Q(\dpath.RF.R[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_110_clk),
    .D(net1977),
    .Q(\dpath.RF.R[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_137_clk),
    .D(net1595),
    .Q(\dpath.RF.R[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_136_clk),
    .D(net2315),
    .Q(\dpath.RF.R[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_111_clk),
    .D(net2191),
    .Q(\dpath.RF.R[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_82_clk),
    .D(net1463),
    .Q(\dpath.RF.R[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_146_clk),
    .D(net1329),
    .Q(\dpath.RF.R[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_81_clk),
    .D(net1799),
    .Q(\dpath.RF.R[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_69_clk),
    .D(net1563),
    .Q(\dpath.RF.R[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_68_clk),
    .D(net1693),
    .Q(\dpath.RF.R[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_72_clk),
    .D(net2337),
    .Q(\dpath.RF.R[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_76_clk),
    .D(net2687),
    .Q(\dpath.RF.R[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_29_clk),
    .D(net1515),
    .Q(\dpath.RF.R[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_26_clk),
    .D(net1405),
    .Q(\dpath.RF.R[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_40_clk),
    .D(net3099),
    .Q(\dpath.RF.R[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_183_clk),
    .D(net1319),
    .Q(\dpath.RF.R[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_180_clk),
    .D(net2077),
    .Q(\dpath.RF.R[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_157_clk),
    .D(net1399),
    .Q(\dpath.RF.R[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_3_clk),
    .D(net2455),
    .Q(\dpath.RF.R[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_176_clk),
    .D(net2935),
    .Q(\dpath.RF.R[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_39_clk),
    .D(net1275),
    .Q(\dpath.RF.R[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_27_clk),
    .D(net2057),
    .Q(\dpath.RF.R[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_36_clk),
    .D(net1717),
    .Q(\dpath.RF.R[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_176_clk),
    .D(net1889),
    .Q(\dpath.RF.R[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_161_clk),
    .D(net1507),
    .Q(\dpath.RF.R[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_172_clk),
    .D(net2169),
    .Q(\dpath.RF.R[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_150_clk),
    .D(net1695),
    .Q(\dpath.RF.R[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_164_clk),
    .D(net1653),
    .Q(\dpath.RF.R[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_123_clk),
    .D(net2717),
    .Q(\dpath.RF.R[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_126_clk),
    .D(net2161),
    .Q(\dpath.RF.R[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_113_clk),
    .D(net1569),
    .Q(\dpath.RF.R[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_127_clk),
    .D(net2107),
    .Q(\dpath.RF.R[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_114_clk),
    .D(net1701),
    .Q(\dpath.RF.R[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_112_clk),
    .D(net1875),
    .Q(\dpath.RF.R[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_142_clk),
    .D(net1489),
    .Q(\dpath.RF.R[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_135_clk),
    .D(net2147),
    .Q(\dpath.RF.R[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_132_clk),
    .D(net1321),
    .Q(\dpath.RF.R[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_133_clk),
    .D(net2207),
    .Q(\dpath.RF.R[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_147_clk),
    .D(net2733),
    .Q(\dpath.RF.R[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_80_clk),
    .D(net2757),
    .Q(\dpath.RF.R[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_69_clk),
    .D(net1495),
    .Q(\dpath.RF.R[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_68_clk),
    .D(net1709),
    .Q(\dpath.RF.R[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_144_clk),
    .D(net2325),
    .Q(\dpath.RF.R[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_76_clk),
    .D(net2891),
    .Q(\dpath.RF.R[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_21_clk),
    .D(net1425),
    .Q(\dpath.RF.R[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_3_clk),
    .D(net1639),
    .Q(\dpath.RF.R[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_29_clk),
    .D(net1197),
    .Q(\dpath.RF.R[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_187_clk),
    .D(net1299),
    .Q(\dpath.RF.R[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_0_clk),
    .D(net2177),
    .Q(\dpath.RF.R[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_178_clk),
    .D(net2483),
    .Q(\dpath.RF.R[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_188_clk),
    .D(net1229),
    .Q(\dpath.RF.R[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_186_clk),
    .D(net1241),
    .Q(\dpath.RF.R[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_33_clk),
    .D(net2027),
    .Q(\dpath.RF.R[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_155_clk),
    .D(net2587),
    .Q(\dpath.RF.R[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_35_clk),
    .D(net1401),
    .Q(\dpath.RF.R[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_175_clk),
    .D(net1713),
    .Q(\dpath.RF.R[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_159_clk),
    .D(net1261),
    .Q(\dpath.RF.R[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_172_clk),
    .D(net2395),
    .Q(\dpath.RF.R[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_153_clk),
    .D(net2181),
    .Q(\dpath.RF.R[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_170_clk),
    .D(net2345),
    .Q(\dpath.RF.R[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_119_clk),
    .D(net2021),
    .Q(\dpath.RF.R[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_168_clk),
    .D(net1533),
    .Q(\dpath.RF.R[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_114_clk),
    .D(net1967),
    .Q(\dpath.RF.R[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_162_clk),
    .D(net1433),
    .Q(\dpath.RF.R[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_116_clk),
    .D(net2767),
    .Q(\dpath.RF.R[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_109_clk),
    .D(net2545),
    .Q(\dpath.RF.R[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_139_clk),
    .D(net1455),
    .Q(\dpath.RF.R[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_128_clk),
    .D(net1231),
    .Q(\dpath.RF.R[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_110_clk),
    .D(net1193),
    .Q(\dpath.RF.R[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_103_clk),
    .D(net1523),
    .Q(\dpath.RF.R[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_148_clk),
    .D(net1857),
    .Q(\dpath.RF.R[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_85_clk),
    .D(net2779),
    .Q(\dpath.RF.R[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_79_clk),
    .D(net1213),
    .Q(\dpath.RF.R[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_77_clk),
    .D(net1427),
    .Q(\dpath.RF.R[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_142_clk),
    .D(net2125),
    .Q(\dpath.RF.R[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_88_clk),
    .D(net2115),
    .Q(\dpath.RF.R[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_20_clk),
    .D(net2159),
    .Q(\dpath.RF.R[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_26_clk),
    .D(net3051),
    .Q(\dpath.RF.R[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_31_clk),
    .D(net1421),
    .Q(\dpath.RF.R[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_180_clk),
    .D(net1491),
    .Q(\dpath.RF.R[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_178_clk),
    .D(net1499),
    .Q(\dpath.RF.R[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_156_clk),
    .D(net1311),
    .Q(\dpath.RF.R[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_25_clk),
    .D(net1233),
    .Q(\dpath.RF.R[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_176_clk),
    .D(net1747),
    .Q(\dpath.RF.R[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_36_clk),
    .D(net1357),
    .Q(\dpath.RF.R[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_154_clk),
    .D(net1395),
    .Q(\dpath.RF.R[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_38_clk),
    .D(net1215),
    .Q(\dpath.RF.R[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_177_clk),
    .D(net1527),
    .Q(\dpath.RF.R[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_162_clk),
    .D(net2005),
    .Q(\dpath.RF.R[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_165_clk),
    .D(net1885),
    .Q(\dpath.RF.R[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_151_clk),
    .D(net2243),
    .Q(\dpath.RF.R[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.CLK(clknet_leaf_166_clk),
    .D(net1359),
    .Q(\dpath.RF.R[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_118_clk),
    .D(net1435),
    .Q(\dpath.RF.R[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_125_clk),
    .D(net2571),
    .Q(\dpath.RF.R[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_114_clk),
    .D(net2515),
    .Q(\dpath.RF.R[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_128_clk),
    .D(net2449),
    .Q(\dpath.RF.R[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_108_clk),
    .D(net1303),
    .Q(\dpath.RF.R[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_110_clk),
    .D(net1279),
    .Q(\dpath.RF.R[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_136_clk),
    .D(net1827),
    .Q(\dpath.RF.R[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_136_clk),
    .D(net2265),
    .Q(\dpath.RF.R[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_111_clk),
    .D(net2457),
    .Q(\dpath.RF.R[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_83_clk),
    .D(net2351),
    .Q(\dpath.RF.R[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_70_clk),
    .D(net3039),
    .Q(\dpath.RF.R[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_84_clk),
    .D(net1631),
    .Q(\dpath.RF.R[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_69_clk),
    .D(net1991),
    .Q(\dpath.RF.R[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_68_clk),
    .D(net1525),
    .Q(\dpath.RF.R[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_72_clk),
    .D(net1553),
    .Q(\dpath.RF.R[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_88_clk),
    .D(net2359),
    .Q(\dpath.RF.R[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_22_clk),
    .D(net3019),
    .Q(\dpath.RF.R[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_3_clk),
    .D(net3037),
    .Q(\dpath.RF.R[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_29_clk),
    .D(net2255),
    .Q(\dpath.RF.R[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_187_clk),
    .D(net2105),
    .Q(\dpath.RF.R[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_0_clk),
    .D(net3033),
    .Q(\dpath.RF.R[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_158_clk),
    .D(net2909),
    .Q(\dpath.RF.R[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_3_clk),
    .D(net2609),
    .Q(\dpath.RF.R[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_185_clk),
    .D(net2881),
    .Q(\dpath.RF.R[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_34_clk),
    .D(net1353),
    .Q(\dpath.RF.R[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_155_clk),
    .D(net2017),
    .Q(\dpath.RF.R[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_149_clk),
    .D(net3035),
    .Q(\dpath.RF.R[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_176_clk),
    .D(net2605),
    .Q(\dpath.RF.R[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_160_clk),
    .D(net2725),
    .Q(\dpath.RF.R[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_171_clk),
    .D(net2489),
    .Q(\dpath.RF.R[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_152_clk),
    .D(net2267),
    .Q(\dpath.RF.R[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_168_clk),
    .D(net2679),
    .Q(\dpath.RF.R[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_123_clk),
    .D(net2947),
    .Q(\dpath.RF.R[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_122_clk),
    .D(net2269),
    .Q(\dpath.RF.R[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_116_clk),
    .D(net3015),
    .Q(\dpath.RF.R[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_125_clk),
    .D(net2109),
    .Q(\dpath.RF.R[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14382_ (.CLK(clknet_leaf_115_clk),
    .D(net3139),
    .Q(\dpath.RF.R[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_110_clk),
    .D(net2859),
    .Q(\dpath.RF.R[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14384_ (.CLK(clknet_leaf_152_clk),
    .D(net2937),
    .Q(\dpath.RF.R[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14385_ (.CLK(clknet_leaf_131_clk),
    .D(net2883),
    .Q(\dpath.RF.R[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14386_ (.CLK(clknet_leaf_111_clk),
    .D(net2871),
    .Q(\dpath.RF.R[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14387_ (.CLK(clknet_leaf_83_clk),
    .D(net2873),
    .Q(\dpath.RF.R[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14388_ (.CLK(clknet_leaf_145_clk),
    .D(net2677),
    .Q(\dpath.RF.R[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_84_clk),
    .D(net2863),
    .Q(\dpath.RF.R[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_73_clk),
    .D(net2431),
    .Q(\dpath.RF.R[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_87_clk),
    .D(net2241),
    .Q(\dpath.RF.R[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_143_clk),
    .D(net2025),
    .Q(\dpath.RF.R[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_88_clk),
    .D(net2175),
    .Q(\dpath.RF.R[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_20_clk),
    .D(net1487),
    .Q(\dpath.RF.R[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_26_clk),
    .D(net1987),
    .Q(\dpath.RF.R[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_31_clk),
    .D(net2221),
    .Q(\dpath.RF.R[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_183_clk),
    .D(net1277),
    .Q(\dpath.RF.R[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_180_clk),
    .D(net1675),
    .Q(\dpath.RF.R[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_156_clk),
    .D(net2187),
    .Q(\dpath.RF.R[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_24_clk),
    .D(net2631),
    .Q(\dpath.RF.R[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_184_clk),
    .D(net1337),
    .Q(\dpath.RF.R[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_33_clk),
    .D(net1305),
    .Q(\dpath.RF.R[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_27_clk),
    .D(net1821),
    .Q(\dpath.RF.R[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_37_clk),
    .D(net1855),
    .Q(\dpath.RF.R[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_177_clk),
    .D(net1677),
    .Q(\dpath.RF.R[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_162_clk),
    .D(net2761),
    .Q(\dpath.RF.R[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_172_clk),
    .D(net1865),
    .Q(\dpath.RF.R[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_151_clk),
    .D(net2729),
    .Q(\dpath.RF.R[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_166_clk),
    .D(net1643),
    .Q(\dpath.RF.R[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.CLK(clknet_leaf_123_clk),
    .D(net2311),
    .Q(\dpath.RF.R[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_122_clk),
    .D(net1873),
    .Q(\dpath.RF.R[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_114_clk),
    .D(net1479),
    .Q(\dpath.RF.R[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_127_clk),
    .D(net1371),
    .Q(\dpath.RF.R[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_114_clk),
    .D(net1539),
    .Q(\dpath.RF.R[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_112_clk),
    .D(net2023),
    .Q(\dpath.RF.R[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_137_clk),
    .D(net1397),
    .Q(\dpath.RF.R[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_136_clk),
    .D(net1737),
    .Q(\dpath.RF.R[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_111_clk),
    .D(net1793),
    .Q(\dpath.RF.R[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_82_clk),
    .D(net1443),
    .Q(\dpath.RF.R[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_147_clk),
    .D(net3109),
    .Q(\dpath.RF.R[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_80_clk),
    .D(net1205),
    .Q(\dpath.RF.R[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_69_clk),
    .D(net1975),
    .Q(\dpath.RF.R[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_68_clk),
    .D(net1385),
    .Q(\dpath.RF.R[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_72_clk),
    .D(net1369),
    .Q(\dpath.RF.R[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_76_clk),
    .D(net1781),
    .Q(\dpath.RF.R[18][31] ));
 sky130_fd_sc_hd__dfxtp_4 _14426_ (.CLK(clknet_leaf_9_clk),
    .D(net3477),
    .Q(net250));
 sky130_fd_sc_hd__dfxtp_2 _14427_ (.CLK(clknet_leaf_9_clk),
    .D(net3494),
    .Q(net253));
 sky130_fd_sc_hd__dfxtp_2 _14428_ (.CLK(clknet_leaf_4_clk),
    .D(net3480),
    .Q(net254));
 sky130_fd_sc_hd__dfxtp_2 _14429_ (.CLK(clknet_leaf_4_clk),
    .D(_00641_),
    .Q(net255));
 sky130_fd_sc_hd__dfxtp_2 _14430_ (.CLK(clknet_leaf_6_clk),
    .D(net3584),
    .Q(net256));
 sky130_fd_sc_hd__dfxtp_2 _14431_ (.CLK(clknet_leaf_6_clk),
    .D(net3515),
    .Q(net257));
 sky130_fd_sc_hd__dfxtp_2 _14432_ (.CLK(clknet_leaf_6_clk),
    .D(net3474),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_6_clk),
    .D(_00645_),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_2 _14434_ (.CLK(clknet_leaf_6_clk),
    .D(net3588),
    .Q(net229));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_6_clk),
    .D(_00647_),
    .Q(net230));
 sky130_fd_sc_hd__dfxtp_2 _14436_ (.CLK(clknet_leaf_7_clk),
    .D(net3580),
    .Q(net231));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_7_clk),
    .D(net3540),
    .Q(net232));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_7_clk),
    .D(net3556),
    .Q(net233));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_7_clk),
    .D(net3511),
    .Q(net234));
 sky130_fd_sc_hd__dfxtp_2 _14440_ (.CLK(clknet_leaf_8_clk),
    .D(net3559),
    .Q(net235));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_8_clk),
    .D(net3545),
    .Q(net236));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_8_clk),
    .D(net3576),
    .Q(net237));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_8_clk),
    .D(net3526),
    .Q(net238));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_11_clk),
    .D(net3538),
    .Q(net240));
 sky130_fd_sc_hd__dfxtp_2 _14445_ (.CLK(clknet_leaf_10_clk),
    .D(net3374),
    .Q(net241));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_11_clk),
    .D(net3398),
    .Q(net242));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_12_clk),
    .D(net3547),
    .Q(net243));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_12_clk),
    .D(net3395),
    .Q(net244));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_10_clk),
    .D(net3508),
    .Q(net245));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_15_clk),
    .D(net3369),
    .Q(net246));
 sky130_fd_sc_hd__dfxtp_2 _14451_ (.CLK(clknet_leaf_15_clk),
    .D(net3254),
    .Q(net247));
 sky130_fd_sc_hd__dfxtp_2 _14452_ (.CLK(clknet_leaf_17_clk),
    .D(net3472),
    .Q(net248));
 sky130_fd_sc_hd__dfxtp_2 _14453_ (.CLK(clknet_leaf_16_clk),
    .D(net3492),
    .Q(net249));
 sky130_fd_sc_hd__dfxtp_2 _14454_ (.CLK(clknet_leaf_18_clk),
    .D(net3225),
    .Q(net251));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_14_clk),
    .D(_00667_),
    .Q(net252));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_20_clk),
    .D(net2097),
    .Q(\dpath.RF.R[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_26_clk),
    .D(net3069),
    .Q(\dpath.RF.R[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_30_clk),
    .D(net3147),
    .Q(\dpath.RF.R[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_182_clk),
    .D(net2877),
    .Q(\dpath.RF.R[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_181_clk),
    .D(net2527),
    .Q(\dpath.RF.R[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_179_clk),
    .D(net2037),
    .Q(\dpath.RF.R[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_3_clk),
    .D(net3137),
    .Q(\dpath.RF.R[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_184_clk),
    .D(net2855),
    .Q(\dpath.RF.R[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_32_clk),
    .D(net2463),
    .Q(\dpath.RF.R[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_26_clk),
    .D(net3005),
    .Q(\dpath.RF.R[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_36_clk),
    .D(net2119),
    .Q(\dpath.RF.R[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_176_clk),
    .D(net3155),
    .Q(\dpath.RF.R[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_161_clk),
    .D(net2699),
    .Q(\dpath.RF.R[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_172_clk),
    .D(net1965),
    .Q(\dpath.RF.R[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_154_clk),
    .D(net2451),
    .Q(\dpath.RF.R[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_165_clk),
    .D(net2053),
    .Q(\dpath.RF.R[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_123_clk),
    .D(net2519),
    .Q(\dpath.RF.R[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_167_clk),
    .D(net1769),
    .Q(\dpath.RF.R[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_130_clk),
    .D(net1483),
    .Q(\dpath.RF.R[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_138_clk),
    .D(net2461),
    .Q(\dpath.RF.R[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_114_clk),
    .D(net2659),
    .Q(\dpath.RF.R[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_113_clk),
    .D(net2673),
    .Q(\dpath.RF.R[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_140_clk),
    .D(net1625),
    .Q(\dpath.RF.R[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_137_clk),
    .D(net3067),
    .Q(\dpath.RF.R[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_131_clk),
    .D(net2823),
    .Q(\dpath.RF.R[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_133_clk),
    .D(net2491),
    .Q(\dpath.RF.R[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_147_clk),
    .D(net3197),
    .Q(\dpath.RF.R[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_79_clk),
    .D(net2409),
    .Q(\dpath.RF.R[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_69_clk),
    .D(net1895),
    .Q(\dpath.RF.R[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_69_clk),
    .D(net2083),
    .Q(\dpath.RF.R[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_146_clk),
    .D(net2289),
    .Q(\dpath.RF.R[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_75_clk),
    .D(net2167),
    .Q(\dpath.RF.R[23][31] ));
 sky130_fd_sc_hd__dfxtp_4 _14488_ (.CLK(clknet_leaf_48_clk),
    .D(_00700_),
    .Q(_00000_));
 sky130_fd_sc_hd__dfxtp_4 _14489_ (.CLK(clknet_leaf_48_clk),
    .D(_00701_),
    .Q(_00001_));
 sky130_fd_sc_hd__dfxtp_4 _14490_ (.CLK(clknet_leaf_46_clk),
    .D(_00702_),
    .Q(_00002_));
 sky130_fd_sc_hd__dfxtp_4 _14491_ (.CLK(clknet_leaf_18_clk),
    .D(_00703_),
    .Q(_00003_));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_17_clk),
    .D(_00704_),
    .Q(_00004_));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_22_clk),
    .D(net1185),
    .Q(\dpath.RF.R[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_24_clk),
    .D(net2963),
    .Q(\dpath.RF.R[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_29_clk),
    .D(net2649),
    .Q(\dpath.RF.R[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_186_clk),
    .D(net1835),
    .Q(\dpath.RF.R[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_0_clk),
    .D(net1379),
    .Q(\dpath.RF.R[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_178_clk),
    .D(net1685),
    .Q(\dpath.RF.R[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_3_clk),
    .D(net2737),
    .Q(\dpath.RF.R[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_185_clk),
    .D(net2919),
    .Q(\dpath.RF.R[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_35_clk),
    .D(net1605),
    .Q(\dpath.RF.R[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_155_clk),
    .D(net2995),
    .Q(\dpath.RF.R[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_150_clk),
    .D(net2271),
    .Q(\dpath.RF.R[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_175_clk),
    .D(net2547),
    .Q(\dpath.RF.R[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_160_clk),
    .D(net1905),
    .Q(\dpath.RF.R[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_173_clk),
    .D(net1621),
    .Q(\dpath.RF.R[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_161_clk),
    .D(net2101),
    .Q(\dpath.RF.R[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_169_clk),
    .D(net1565),
    .Q(\dpath.RF.R[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_119_clk),
    .D(net2309),
    .Q(\dpath.RF.R[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_120_clk),
    .D(net2667),
    .Q(\dpath.RF.R[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_116_clk),
    .D(net2343),
    .Q(\dpath.RF.R[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_126_clk),
    .D(net1445),
    .Q(\dpath.RF.R[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_116_clk),
    .D(net3003),
    .Q(\dpath.RF.R[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_109_clk),
    .D(net2379),
    .Q(\dpath.RF.R[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_162_clk),
    .D(net2121),
    .Q(\dpath.RF.R[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_131_clk),
    .D(net1545),
    .Q(\dpath.RF.R[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_103_clk),
    .D(net2807),
    .Q(\dpath.RF.R[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_102_clk),
    .D(net1327),
    .Q(\dpath.RF.R[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_140_clk),
    .D(net1579),
    .Q(\dpath.RF.R[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_85_clk),
    .D(net1745),
    .Q(\dpath.RF.R[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_78_clk),
    .D(net1245),
    .Q(\dpath.RF.R[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_87_clk),
    .D(net1309),
    .Q(\dpath.RF.R[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_136_clk),
    .D(net1771),
    .Q(\dpath.RF.R[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_89_clk),
    .D(net1281),
    .Q(\dpath.RF.R[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_21_clk),
    .D(net1335),
    .Q(\dpath.RF.R[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_25_clk),
    .D(net2885),
    .Q(\dpath.RF.R[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_30_clk),
    .D(net1375),
    .Q(\dpath.RF.R[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_181_clk),
    .D(net3059),
    .Q(\dpath.RF.R[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_1_clk),
    .D(net3091),
    .Q(\dpath.RF.R[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_158_clk),
    .D(net3135),
    .Q(\dpath.RF.R[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_2_clk),
    .D(net2903),
    .Q(\dpath.RF.R[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_182_clk),
    .D(net1797),
    .Q(\dpath.RF.R[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_33_clk),
    .D(net2681),
    .Q(\dpath.RF.R[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_27_clk),
    .D(net1645),
    .Q(\dpath.RF.R[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_35_clk),
    .D(net2879),
    .Q(\dpath.RF.R[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_178_clk),
    .D(net3073),
    .Q(\dpath.RF.R[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_160_clk),
    .D(net3161),
    .Q(\dpath.RF.R[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_177_clk),
    .D(net2397),
    .Q(\dpath.RF.R[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_153_clk),
    .D(net1549),
    .Q(\dpath.RF.R[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_165_clk),
    .D(net2469),
    .Q(\dpath.RF.R[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_125_clk),
    .D(net2819),
    .Q(\dpath.RF.R[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_163_clk),
    .D(net1589),
    .Q(\dpath.RF.R[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_129_clk),
    .D(net1963),
    .Q(\dpath.RF.R[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_126_clk),
    .D(net2529),
    .Q(\dpath.RF.R[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_113_clk),
    .D(net2357),
    .Q(\dpath.RF.R[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_113_clk),
    .D(net2307),
    .Q(\dpath.RF.R[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_138_clk),
    .D(net2773),
    .Q(\dpath.RF.R[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_134_clk),
    .D(net2383),
    .Q(\dpath.RF.R[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_132_clk),
    .D(net2045),
    .Q(\dpath.RF.R[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_133_clk),
    .D(net1879),
    .Q(\dpath.RF.R[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_148_clk),
    .D(net1723),
    .Q(\dpath.RF.R[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_80_clk),
    .D(net1765),
    .Q(\dpath.RF.R[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_75_clk),
    .D(net2387),
    .Q(\dpath.RF.R[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_76_clk),
    .D(net3095),
    .Q(\dpath.RF.R[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_144_clk),
    .D(net2791),
    .Q(\dpath.RF.R[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_78_clk),
    .D(net2537),
    .Q(\dpath.RF.R[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_21_clk),
    .D(net1061),
    .Q(\dpath.RF.R[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_3_clk),
    .D(net1147),
    .Q(\dpath.RF.R[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_30_clk),
    .D(net1171),
    .Q(\dpath.RF.R[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_187_clk),
    .D(net1099),
    .Q(\dpath.RF.R[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_0_clk),
    .D(net1081),
    .Q(\dpath.RF.R[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_178_clk),
    .D(net1159),
    .Q(\dpath.RF.R[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_188_clk),
    .D(net1083),
    .Q(\dpath.RF.R[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_186_clk),
    .D(net1075),
    .Q(\dpath.RF.R[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_33_clk),
    .D(net1115),
    .Q(\dpath.RF.R[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_155_clk),
    .D(net1121),
    .Q(\dpath.RF.R[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_149_clk),
    .D(net1125),
    .Q(\dpath.RF.R[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_175_clk),
    .D(net1149),
    .Q(\dpath.RF.R[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_159_clk),
    .D(net1143),
    .Q(\dpath.RF.R[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_172_clk),
    .D(net1131),
    .Q(\dpath.RF.R[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_152_clk),
    .D(net1127),
    .Q(\dpath.RF.R[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_170_clk),
    .D(net1145),
    .Q(\dpath.RF.R[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_120_clk),
    .D(net1179),
    .Q(\dpath.RF.R[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_168_clk),
    .D(net1119),
    .Q(\dpath.RF.R[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_114_clk),
    .D(net1135),
    .Q(\dpath.RF.R[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_126_clk),
    .D(net1113),
    .Q(\dpath.RF.R[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_116_clk),
    .D(net1103),
    .Q(\dpath.RF.R[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_109_clk),
    .D(net1097),
    .Q(\dpath.RF.R[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_139_clk),
    .D(net1101),
    .Q(\dpath.RF.R[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_131_clk),
    .D(net1165),
    .Q(\dpath.RF.R[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_4_11__leaf_clk),
    .D(net1175),
    .Q(\dpath.RF.R[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_102_clk),
    .D(net1059),
    .Q(\dpath.RF.R[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_148_clk),
    .D(net1137),
    .Q(\dpath.RF.R[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_85_clk),
    .D(net1053),
    .Q(\dpath.RF.R[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_78_clk),
    .D(net1155),
    .Q(\dpath.RF.R[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_77_clk),
    .D(net1161),
    .Q(\dpath.RF.R[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_142_clk),
    .D(net1109),
    .Q(\dpath.RF.R[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_88_clk),
    .D(net1123),
    .Q(\dpath.RF.R[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_16_clk),
    .D(net2787),
    .Q(\dpath.RF.R[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_4_clk),
    .D(net1803),
    .Q(\dpath.RF.R[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_20_clk),
    .D(net2297),
    .Q(\dpath.RF.R[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_187_clk),
    .D(net1867),
    .Q(\dpath.RF.R[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_188_clk),
    .D(net1757),
    .Q(\dpath.RF.R[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_178_clk),
    .D(net2237),
    .Q(\dpath.RF.R[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_188_clk),
    .D(net2845),
    .Q(\dpath.RF.R[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_186_clk),
    .D(net2441),
    .Q(\dpath.RF.R[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_33_clk),
    .D(net2213),
    .Q(\dpath.RF.R[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_156_clk),
    .D(net2475),
    .Q(\dpath.RF.R[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_35_clk),
    .D(net2087),
    .Q(\dpath.RF.R[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_175_clk),
    .D(net2085),
    .Q(\dpath.RF.R[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_158_clk),
    .D(net2091),
    .Q(\dpath.RF.R[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_172_clk),
    .D(net1593),
    .Q(\dpath.RF.R[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_153_clk),
    .D(net2485),
    .Q(\dpath.RF.R[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_171_clk),
    .D(net2333),
    .Q(\dpath.RF.R[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_122_clk),
    .D(net1481),
    .Q(\dpath.RF.R[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_168_clk),
    .D(net2293),
    .Q(\dpath.RF.R[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_118_clk),
    .D(net1437),
    .Q(\dpath.RF.R[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_162_clk),
    .D(net1509),
    .Q(\dpath.RF.R[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_116_clk),
    .D(net2805),
    .Q(\dpath.RF.R[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_109_clk),
    .D(net2401),
    .Q(\dpath.RF.R[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_139_clk),
    .D(net1403),
    .Q(\dpath.RF.R[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_128_clk),
    .D(net2019),
    .Q(\dpath.RF.R[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_110_clk),
    .D(net1207),
    .Q(\dpath.RF.R[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_103_clk),
    .D(net1381),
    .Q(\dpath.RF.R[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_150_clk),
    .D(net2141),
    .Q(\dpath.RF.R[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_84_clk),
    .D(net1519),
    .Q(\dpath.RF.R[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_143_clk),
    .D(net1599),
    .Q(\dpath.RF.R[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_78_clk),
    .D(net1929),
    .Q(\dpath.RF.R[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_140_clk),
    .D(net1249),
    .Q(\dpath.RF.R[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_88_clk),
    .D(net1453),
    .Q(\dpath.RF.R[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_22_clk),
    .D(net1751),
    .Q(\dpath.RF.R[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_24_clk),
    .D(net2851),
    .Q(\dpath.RF.R[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_27_clk),
    .D(net1659),
    .Q(\dpath.RF.R[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_186_clk),
    .D(net1819),
    .Q(\dpath.RF.R[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_0_clk),
    .D(net1417),
    .Q(\dpath.RF.R[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_178_clk),
    .D(net2389),
    .Q(\dpath.RF.R[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_4_clk),
    .D(net1891),
    .Q(\dpath.RF.R[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_185_clk),
    .D(net2411),
    .Q(\dpath.RF.R[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_28_clk),
    .D(net1271),
    .Q(\dpath.RF.R[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_155_clk),
    .D(net1465),
    .Q(\dpath.RF.R[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_149_clk),
    .D(net1953),
    .Q(\dpath.RF.R[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_175_clk),
    .D(net2593),
    .Q(\dpath.RF.R[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_160_clk),
    .D(net2123),
    .Q(\dpath.RF.R[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_173_clk),
    .D(net2047),
    .Q(\dpath.RF.R[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_161_clk),
    .D(net1783),
    .Q(\dpath.RF.R[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_170_clk),
    .D(net2581),
    .Q(\dpath.RF.R[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_119_clk),
    .D(net2279),
    .Q(\dpath.RF.R[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_121_clk),
    .D(net1247),
    .Q(\dpath.RF.R[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_117_clk),
    .D(net2153),
    .Q(\dpath.RF.R[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_126_clk),
    .D(net2453),
    .Q(\dpath.RF.R[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_116_clk),
    .D(net1511),
    .Q(\dpath.RF.R[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_108_clk),
    .D(net1219),
    .Q(\dpath.RF.R[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_162_clk),
    .D(net2961),
    .Q(\dpath.RF.R[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_131_clk),
    .D(net1743),
    .Q(\dpath.RF.R[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_111_clk),
    .D(net1815),
    .Q(\dpath.RF.R[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_83_clk),
    .D(net1191),
    .Q(\dpath.RF.R[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_151_clk),
    .D(net2705),
    .Q(\dpath.RF.R[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_84_clk),
    .D(net1377),
    .Q(\dpath.RF.R[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_78_clk),
    .D(net1259),
    .Q(\dpath.RF.R[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_87_clk),
    .D(net1623),
    .Q(\dpath.RF.R[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_142_clk),
    .D(net1237),
    .Q(\dpath.RF.R[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_87_clk),
    .D(net1683),
    .Q(\dpath.RF.R[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_23_clk),
    .D(net3085),
    .Q(\dpath.RF.R[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_26_clk),
    .D(net1749),
    .Q(\dpath.RF.R[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_33_clk),
    .D(net1349),
    .Q(\dpath.RF.R[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_180_clk),
    .D(net1853),
    .Q(\dpath.RF.R[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_179_clk),
    .D(net2513),
    .Q(\dpath.RF.R[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_158_clk),
    .D(net1331),
    .Q(\dpath.RF.R[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_179_clk),
    .D(net1361),
    .Q(\dpath.RF.R[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_178_clk),
    .D(net1995),
    .Q(\dpath.RF.R[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_33_clk),
    .D(net2683),
    .Q(\dpath.RF.R[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_154_clk),
    .D(net2199),
    .Q(\dpath.RF.R[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_147_clk),
    .D(net1861),
    .Q(\dpath.RF.R[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_177_clk),
    .D(net2145),
    .Q(\dpath.RF.R[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_162_clk),
    .D(net1893),
    .Q(\dpath.RF.R[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_165_clk),
    .D(net1493),
    .Q(\dpath.RF.R[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_152_clk),
    .D(net1687),
    .Q(\dpath.RF.R[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_163_clk),
    .D(net2143),
    .Q(\dpath.RF.R[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_130_clk),
    .D(net2327),
    .Q(\dpath.RF.R[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_125_clk),
    .D(net1955),
    .Q(\dpath.RF.R[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_131_clk),
    .D(net2231),
    .Q(\dpath.RF.R[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_129_clk),
    .D(net1617),
    .Q(\dpath.RF.R[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_112_clk),
    .D(net2089),
    .Q(\dpath.RF.R[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_110_clk),
    .D(net1817),
    .Q(\dpath.RF.R[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_137_clk),
    .D(net1341),
    .Q(\dpath.RF.R[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_135_clk),
    .D(net1503),
    .Q(\dpath.RF.R[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_111_clk),
    .D(net1667),
    .Q(\dpath.RF.R[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_133_clk),
    .D(net1973),
    .Q(\dpath.RF.R[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_145_clk),
    .D(net2569),
    .Q(\dpath.RF.R[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_81_clk),
    .D(net2669),
    .Q(\dpath.RF.R[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_74_clk),
    .D(net1547),
    .Q(\dpath.RF.R[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_88_clk),
    .D(net1773),
    .Q(\dpath.RF.R[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_72_clk),
    .D(net1383),
    .Q(\dpath.RF.R[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_77_clk),
    .D(net1365),
    .Q(\dpath.RF.R[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_17_clk),
    .D(net2275),
    .Q(\dpath.RF.R[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_25_clk),
    .D(net1239),
    .Q(\dpath.RF.R[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_30_clk),
    .D(net2149),
    .Q(\dpath.RF.R[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_181_clk),
    .D(net1615),
    .Q(\dpath.RF.R[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_1_clk),
    .D(net1567),
    .Q(\dpath.RF.R[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_179_clk),
    .D(net2111),
    .Q(\dpath.RF.R[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_1_clk),
    .D(net2185),
    .Q(\dpath.RF.R[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_181_clk),
    .D(net1439),
    .Q(\dpath.RF.R[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_32_clk),
    .D(net1711),
    .Q(\dpath.RF.R[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_27_clk),
    .D(net1475),
    .Q(\dpath.RF.R[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_36_clk),
    .D(net1325),
    .Q(\dpath.RF.R[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_178_clk),
    .D(net2281),
    .Q(\dpath.RF.R[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_160_clk),
    .D(net2811),
    .Q(\dpath.RF.R[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_177_clk),
    .D(net2651),
    .Q(\dpath.RF.R[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_153_clk),
    .D(net1911),
    .Q(\dpath.RF.R[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_165_clk),
    .D(net1633),
    .Q(\dpath.RF.R[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_125_clk),
    .D(net1883),
    .Q(\dpath.RF.R[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_163_clk),
    .D(net2435),
    .Q(\dpath.RF.R[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_129_clk),
    .D(net1807),
    .Q(\dpath.RF.R[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_127_clk),
    .D(net1937),
    .Q(\dpath.RF.R[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_114_clk),
    .D(net1829),
    .Q(\dpath.RF.R[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_113_clk),
    .D(net2139),
    .Q(\dpath.RF.R[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_138_clk),
    .D(net1387),
    .Q(\dpath.RF.R[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_135_clk),
    .D(net1221),
    .Q(\dpath.RF.R[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_131_clk),
    .D(net2163),
    .Q(\dpath.RF.R[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_134_clk),
    .D(net1227),
    .Q(\dpath.RF.R[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_148_clk),
    .D(net2429),
    .Q(\dpath.RF.R[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_80_clk),
    .D(net1933),
    .Q(\dpath.RF.R[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_74_clk),
    .D(net1627),
    .Q(\dpath.RF.R[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_75_clk),
    .D(net1409),
    .Q(\dpath.RF.R[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_144_clk),
    .D(net1551),
    .Q(\dpath.RF.R[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_74_clk),
    .D(net1467),
    .Q(\dpath.RF.R[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_22_clk),
    .D(net2499),
    .Q(\dpath.RF.R[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_24_clk),
    .D(net3093),
    .Q(\dpath.RF.R[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_27_clk),
    .D(net2913),
    .Q(\dpath.RF.R[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_186_clk),
    .D(net3115),
    .Q(\dpath.RF.R[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_0_clk),
    .D(net2295),
    .Q(\dpath.RF.R[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_178_clk),
    .D(net2249),
    .Q(\dpath.RF.R[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_6_clk),
    .D(net2889),
    .Q(\dpath.RF.R[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_185_clk),
    .D(net2373),
    .Q(\dpath.RF.R[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_28_clk),
    .D(net1947),
    .Q(\dpath.RF.R[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_155_clk),
    .D(net2481),
    .Q(\dpath.RF.R[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_150_clk),
    .D(net1863),
    .Q(\dpath.RF.R[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_175_clk),
    .D(net3159),
    .Q(\dpath.RF.R[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.CLK(clknet_leaf_160_clk),
    .D(net2983),
    .Q(\dpath.RF.R[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_173_clk),
    .D(net2013),
    .Q(\dpath.RF.R[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_161_clk),
    .D(net2531),
    .Q(\dpath.RF.R[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_170_clk),
    .D(net2303),
    .Q(\dpath.RF.R[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_119_clk),
    .D(net3097),
    .Q(\dpath.RF.R[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_121_clk),
    .D(net2813),
    .Q(\dpath.RF.R[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_117_clk),
    .D(net2943),
    .Q(\dpath.RF.R[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_126_clk),
    .D(net2847),
    .Q(\dpath.RF.R[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_108_clk),
    .D(net2633),
    .Q(\dpath.RF.R[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_108_clk),
    .D(net1761),
    .Q(\dpath.RF.R[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_162_clk),
    .D(net2957),
    .Q(\dpath.RF.R[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.CLK(clknet_leaf_131_clk),
    .D(net3025),
    .Q(\dpath.RF.R[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_103_clk),
    .D(net2137),
    .Q(\dpath.RF.R[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_102_clk),
    .D(net2793),
    .Q(\dpath.RF.R[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_150_clk),
    .D(net2799),
    .Q(\dpath.RF.R[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_85_clk),
    .D(net2001),
    .Q(\dpath.RF.R[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_78_clk),
    .D(net2905),
    .Q(\dpath.RF.R[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_87_clk),
    .D(net1983),
    .Q(\dpath.RF.R[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_136_clk),
    .D(net3165),
    .Q(\dpath.RF.R[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.CLK(clknet_leaf_87_clk),
    .D(net1887),
    .Q(\dpath.RF.R[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_17_clk),
    .D(net3149),
    .Q(\dpath.RF.R[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_25_clk),
    .D(net1901),
    .Q(\dpath.RF.R[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.CLK(clknet_leaf_30_clk),
    .D(net2075),
    .Q(\dpath.RF.R[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14752_ (.CLK(clknet_leaf_181_clk),
    .D(net2205),
    .Q(\dpath.RF.R[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.CLK(clknet_leaf_1_clk),
    .D(net2777),
    .Q(\dpath.RF.R[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.CLK(clknet_leaf_179_clk),
    .D(net2063),
    .Q(\dpath.RF.R[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.CLK(clknet_leaf_1_clk),
    .D(net2341),
    .Q(\dpath.RF.R[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.CLK(clknet_leaf_182_clk),
    .D(net2691),
    .Q(\dpath.RF.R[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.CLK(clknet_leaf_32_clk),
    .D(net2033),
    .Q(\dpath.RF.R[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.CLK(clknet_leaf_27_clk),
    .D(net2417),
    .Q(\dpath.RF.R[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.CLK(clknet_leaf_35_clk),
    .D(net1079),
    .Q(\dpath.RF.R[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.CLK(clknet_leaf_178_clk),
    .D(net3023),
    .Q(\dpath.RF.R[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_160_clk),
    .D(net2857),
    .Q(\dpath.RF.R[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.CLK(clknet_leaf_177_clk),
    .D(net3111),
    .Q(\dpath.RF.R[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_153_clk),
    .D(net2193),
    .Q(\dpath.RF.R[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_165_clk),
    .D(net2695),
    .Q(\dpath.RF.R[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_125_clk),
    .D(net2055),
    .Q(\dpath.RF.R[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_163_clk),
    .D(net2997),
    .Q(\dpath.RF.R[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_129_clk),
    .D(net1759),
    .Q(\dpath.RF.R[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_162_clk),
    .D(net3163),
    .Q(\dpath.RF.R[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_113_clk),
    .D(net2069),
    .Q(\dpath.RF.R[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_113_clk),
    .D(net2335),
    .Q(\dpath.RF.R[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_138_clk),
    .D(net2259),
    .Q(\dpath.RF.R[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_135_clk),
    .D(net2611),
    .Q(\dpath.RF.R[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_131_clk),
    .D(net3143),
    .Q(\dpath.RF.R[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_134_clk),
    .D(net3055),
    .Q(\dpath.RF.R[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.CLK(clknet_leaf_147_clk),
    .D(net2931),
    .Q(\dpath.RF.R[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_80_clk),
    .D(net1669),
    .Q(\dpath.RF.R[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_75_clk),
    .D(net2525),
    .Q(\dpath.RF.R[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_75_clk),
    .D(net2113),
    .Q(\dpath.RF.R[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_144_clk),
    .D(net1691),
    .Q(\dpath.RF.R[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_74_clk),
    .D(net2285),
    .Q(\dpath.RF.R[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_22_clk),
    .D(net1485),
    .Q(\dpath.RF.R[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.CLK(clknet_leaf_23_clk),
    .D(net2693),
    .Q(\dpath.RF.R[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_28_clk),
    .D(net2841),
    .Q(\dpath.RF.R[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_186_clk),
    .D(net1999),
    .Q(\dpath.RF.R[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_181_clk),
    .D(net2471),
    .Q(\dpath.RF.R[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_160_clk),
    .D(net2247),
    .Q(\dpath.RF.R[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_4_clk),
    .D(net1949),
    .Q(\dpath.RF.R[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_185_clk),
    .D(net2835),
    .Q(\dpath.RF.R[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_149_clk),
    .D(net2367),
    .Q(\dpath.RF.R[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_155_clk),
    .D(net1561),
    .Q(\dpath.RF.R[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_150_clk),
    .D(net2479),
    .Q(\dpath.RF.R[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_174_clk),
    .D(net2501),
    .Q(\dpath.RF.R[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_160_clk),
    .D(net2273),
    .Q(\dpath.RF.R[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_171_clk),
    .D(net1681),
    .Q(\dpath.RF.R[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_152_clk),
    .D(net1535),
    .Q(\dpath.RF.R[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_168_clk),
    .D(net1833),
    .Q(\dpath.RF.R[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_118_clk),
    .D(net2477),
    .Q(\dpath.RF.R[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_120_clk),
    .D(net2203),
    .Q(\dpath.RF.R[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_116_clk),
    .D(net2007),
    .Q(\dpath.RF.R[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_125_clk),
    .D(net1351),
    .Q(\dpath.RF.R[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_108_clk),
    .D(net1981),
    .Q(\dpath.RF.R[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_109_clk),
    .D(net2473),
    .Q(\dpath.RF.R[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_139_clk),
    .D(net1689),
    .Q(\dpath.RF.R[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_131_clk),
    .D(net2127),
    .Q(\dpath.RF.R[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_103_clk),
    .D(net2753),
    .Q(\dpath.RF.R[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.CLK(clknet_leaf_102_clk),
    .D(net1195),
    .Q(\dpath.RF.R[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_140_clk),
    .D(net2081),
    .Q(\dpath.RF.R[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_85_clk),
    .D(net1459),
    .Q(\dpath.RF.R[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.CLK(clknet_leaf_78_clk),
    .D(net1267),
    .Q(\dpath.RF.R[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.CLK(clknet_leaf_86_clk),
    .D(net1183),
    .Q(\dpath.RF.R[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_136_clk),
    .D(net3133),
    .Q(\dpath.RF.R[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.CLK(clknet_leaf_89_clk),
    .D(net1265),
    .Q(\dpath.RF.R[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_62_clk),
    .D(_01025_),
    .Q(net324));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.CLK(clknet_leaf_62_clk),
    .D(_01026_),
    .Q(net335));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.CLK(clknet_leaf_63_clk),
    .D(_01027_),
    .Q(net346));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_62_clk),
    .D(_01028_),
    .Q(net349));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.CLK(clknet_leaf_61_clk),
    .D(_01029_),
    .Q(net350));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_62_clk),
    .D(_01030_),
    .Q(net351));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_61_clk),
    .D(_01031_),
    .Q(net352));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_61_clk),
    .D(_01032_),
    .Q(net353));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_61_clk),
    .D(_01033_),
    .Q(net354));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_61_clk),
    .D(_01034_),
    .Q(net355));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_61_clk),
    .D(_01035_),
    .Q(net325));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_61_clk),
    .D(_01036_),
    .Q(net326));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_60_clk),
    .D(_01037_),
    .Q(net327));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_62_clk),
    .D(_01038_),
    .Q(net328));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_62_clk),
    .D(_01039_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_2 _14828_ (.CLK(clknet_leaf_63_clk),
    .D(_01040_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_2 _14829_ (.CLK(clknet_leaf_64_clk),
    .D(_01041_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_2 _14830_ (.CLK(clknet_leaf_64_clk),
    .D(_01042_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_2 _14831_ (.CLK(clknet_leaf_63_clk),
    .D(_01043_),
    .Q(net333));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_61_clk),
    .D(_01044_),
    .Q(net334));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_60_clk),
    .D(_01045_),
    .Q(net336));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_60_clk),
    .D(_01046_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.CLK(clknet_leaf_60_clk),
    .D(_01047_),
    .Q(net338));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_60_clk),
    .D(_01048_),
    .Q(net339));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_60_clk),
    .D(_01049_),
    .Q(net340));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_60_clk),
    .D(_01050_),
    .Q(net341));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_60_clk),
    .D(_01051_),
    .Q(net342));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_61_clk),
    .D(_01052_),
    .Q(net343));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_60_clk),
    .D(_01053_),
    .Q(net344));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_60_clk),
    .D(_01054_),
    .Q(net345));
 sky130_fd_sc_hd__dfxtp_2 _14843_ (.CLK(clknet_leaf_62_clk),
    .D(_01055_),
    .Q(net347));
 sky130_fd_sc_hd__dfxtp_2 _14844_ (.CLK(clknet_leaf_62_clk),
    .D(_01056_),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.CLK(clknet_leaf_94_clk),
    .D(net3383),
    .Q(net292));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.CLK(clknet_leaf_97_clk),
    .D(net3407),
    .Q(net303));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.CLK(clknet_leaf_94_clk),
    .D(net3377),
    .Q(net314));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_94_clk),
    .D(net3409),
    .Q(net317));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_93_clk),
    .D(net3348),
    .Q(net318));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.CLK(clknet_leaf_93_clk),
    .D(net3391),
    .Q(net319));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.CLK(clknet_leaf_93_clk),
    .D(net3329),
    .Q(net320));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_leaf_93_clk),
    .D(net3344),
    .Q(net321));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.CLK(clknet_leaf_93_clk),
    .D(net3331),
    .Q(net322));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.CLK(clknet_leaf_92_clk),
    .D(net3365),
    .Q(net323));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.CLK(clknet_leaf_92_clk),
    .D(net3353),
    .Q(net293));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_92_clk),
    .D(net3320),
    .Q(net294));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_92_clk),
    .D(net3318),
    .Q(net295));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_92_clk),
    .D(net3316),
    .Q(net296));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_92_clk),
    .D(net3314),
    .Q(net297));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_65_clk),
    .D(net3294),
    .Q(net298));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_65_clk),
    .D(net3300),
    .Q(net299));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_64_clk),
    .D(net3333),
    .Q(net300));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_64_clk),
    .D(net3304),
    .Q(net301));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_64_clk),
    .D(net3322),
    .Q(net302));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_64_clk),
    .D(net3371),
    .Q(net304));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_64_clk),
    .D(net3351),
    .Q(net305));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_63_clk),
    .D(net3361),
    .Q(net306));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_63_clk),
    .D(net3363),
    .Q(net307));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_63_clk),
    .D(net3355),
    .Q(net308));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_63_clk),
    .D(net3357),
    .Q(net309));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_63_clk),
    .D(net3389),
    .Q(net310));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_63_clk),
    .D(net3387),
    .Q(net311));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_63_clk),
    .D(net3385),
    .Q(net312));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_63_clk),
    .D(net3414),
    .Q(net313));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_63_clk),
    .D(net3379),
    .Q(net315));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_63_clk),
    .D(net3419),
    .Q(net316));
 sky130_fd_sc_hd__dfxtp_2 _14877_ (.CLK(clknet_leaf_96_clk),
    .D(net3215),
    .Q(net260));
 sky130_fd_sc_hd__dfxtp_2 _14878_ (.CLK(clknet_leaf_97_clk),
    .D(net3258),
    .Q(net271));
 sky130_fd_sc_hd__dfxtp_2 _14879_ (.CLK(clknet_leaf_98_clk),
    .D(net3444),
    .Q(net282));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_106_clk),
    .D(net3482),
    .Q(net285));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_107_clk),
    .D(net3524),
    .Q(net286));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_107_clk),
    .D(net3517),
    .Q(net287));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_107_clk),
    .D(net3549),
    .Q(net288));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_107_clk),
    .D(net3530),
    .Q(net289));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_106_clk),
    .D(net3498),
    .Q(net290));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_106_clk),
    .D(net3503),
    .Q(net291));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_107_clk),
    .D(net3513),
    .Q(net261));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_107_clk),
    .D(net3521),
    .Q(net262));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_107_clk),
    .D(net3533),
    .Q(net263));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_98_clk),
    .D(net3434),
    .Q(net264));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_106_clk),
    .D(net3458),
    .Q(net265));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_106_clk),
    .D(net3405),
    .Q(net266));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_106_clk),
    .D(net3367),
    .Q(net267));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_106_clk),
    .D(net3335),
    .Q(net268));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_106_clk),
    .D(net3248),
    .Q(net269));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_106_clk),
    .D(net3489),
    .Q(net270));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_99_clk),
    .D(net3487),
    .Q(net272));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_99_clk),
    .D(net3501),
    .Q(net273));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_98_clk),
    .D(net3449),
    .Q(net274));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_98_clk),
    .D(net3256),
    .Q(net275));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_98_clk),
    .D(net3218),
    .Q(net276));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_98_clk),
    .D(net3451),
    .Q(net277));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.CLK(clknet_leaf_98_clk),
    .D(net3431),
    .Q(net278));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_97_clk),
    .D(net3381),
    .Q(net279));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_97_clk),
    .D(net3460),
    .Q(net280));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_97_clk),
    .D(net3438),
    .Q(net281));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.CLK(clknet_leaf_97_clk),
    .D(net3506),
    .Q(net283));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_97_clk),
    .D(net3290),
    .Q(net284));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.CLK(clknet_leaf_68_clk),
    .D(_01121_),
    .Q(\dpath.csrw_out_DX.q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_70_clk),
    .D(_01122_),
    .Q(\dpath.csrw_out_DX.q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_148_clk),
    .D(_01123_),
    .Q(\dpath.csrw_out_DX.q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_157_clk),
    .D(_01124_),
    .Q(\dpath.csrw_out_DX.q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_156_clk),
    .D(_01125_),
    .Q(\dpath.csrw_out_DX.q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_153_clk),
    .D(_01126_),
    .Q(\dpath.csrw_out_DX.q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_156_clk),
    .D(_01127_),
    .Q(\dpath.csrw_out_DX.q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_149_clk),
    .D(_01128_),
    .Q(\dpath.csrw_out_DX.q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_85_clk),
    .D(_01129_),
    .Q(\dpath.csrw_out_DX.q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_136_clk),
    .D(_01130_),
    .Q(\dpath.csrw_out_DX.q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_101_clk),
    .D(_01131_),
    .Q(\dpath.csrw_out_DX.q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_153_clk),
    .D(_01132_),
    .Q(\dpath.csrw_out_DX.q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_102_clk),
    .D(_01133_),
    .Q(\dpath.csrw_out_DX.q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_102_clk),
    .D(_01134_),
    .Q(\dpath.csrw_out_DX.q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.CLK(clknet_leaf_100_clk),
    .D(_01135_),
    .Q(\dpath.csrw_out_DX.q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_101_clk),
    .D(_01136_),
    .Q(\dpath.csrw_out_DX.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_105_clk),
    .D(_01137_),
    .Q(\dpath.csrw_out_DX.q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_85_clk),
    .D(_01138_),
    .Q(\dpath.csrw_out_DX.q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14927_ (.CLK(clknet_leaf_105_clk),
    .D(_01139_),
    .Q(\dpath.csrw_out_DX.q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.CLK(clknet_leaf_95_clk),
    .D(_01140_),
    .Q(\dpath.csrw_out_DX.q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14929_ (.CLK(clknet_leaf_100_clk),
    .D(_01141_),
    .Q(\dpath.csrw_out_DX.q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.CLK(clknet_leaf_100_clk),
    .D(_01142_),
    .Q(\dpath.csrw_out_DX.q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_101_clk),
    .D(_01143_),
    .Q(\dpath.csrw_out_DX.q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_91_clk),
    .D(_01144_),
    .Q(\dpath.csrw_out_DX.q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_90_clk),
    .D(_01145_),
    .Q(\dpath.csrw_out_DX.q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_90_clk),
    .D(_01146_),
    .Q(\dpath.csrw_out_DX.q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_90_clk),
    .D(_01147_),
    .Q(\dpath.csrw_out_DX.q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_90_clk),
    .D(_01148_),
    .Q(\dpath.csrw_out_DX.q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_89_clk),
    .D(_01149_),
    .Q(\dpath.csrw_out_DX.q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_71_clk),
    .D(_01150_),
    .Q(\dpath.csrw_out_DX.q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_89_clk),
    .D(_01151_),
    .Q(\dpath.csrw_out_DX.q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_88_clk),
    .D(_01152_),
    .Q(\dpath.csrw_out_DX.q[31] ));
 sky130_fd_sc_hd__dfxtp_4 _14941_ (.CLK(clknet_leaf_44_clk),
    .D(_01153_),
    .Q(\dpath.alu.adder.in1[0] ));
 sky130_fd_sc_hd__dfxtp_4 _14942_ (.CLK(clknet_leaf_43_clk),
    .D(_01154_),
    .Q(\dpath.alu.adder.in1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_31_clk),
    .D(_01155_),
    .Q(\dpath.alu.adder.in1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14944_ (.CLK(clknet_leaf_43_clk),
    .D(_01156_),
    .Q(\dpath.alu.adder.in1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_44_clk),
    .D(_01157_),
    .Q(\dpath.alu.adder.in1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_41_clk),
    .D(_01158_),
    .Q(\dpath.alu.adder.in1[5] ));
 sky130_fd_sc_hd__dfxtp_4 _14947_ (.CLK(clknet_leaf_43_clk),
    .D(_01159_),
    .Q(\dpath.alu.adder.in1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_41_clk),
    .D(_01160_),
    .Q(\dpath.alu.adder.in1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_40_clk),
    .D(_01161_),
    .Q(\dpath.alu.adder.in1[8] ));
 sky130_fd_sc_hd__dfxtp_4 _14950_ (.CLK(clknet_leaf_40_clk),
    .D(_01162_),
    .Q(\dpath.alu.adder.in1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_40_clk),
    .D(_01163_),
    .Q(\dpath.alu.adder.in1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_40_clk),
    .D(_01164_),
    .Q(\dpath.alu.adder.in1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14953_ (.CLK(clknet_leaf_39_clk),
    .D(_01165_),
    .Q(\dpath.alu.adder.in1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14954_ (.CLK(clknet_leaf_39_clk),
    .D(_01166_),
    .Q(\dpath.alu.adder.in1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_37_clk),
    .D(_01167_),
    .Q(\dpath.alu.adder.in1[14] ));
 sky130_fd_sc_hd__dfxtp_4 _14956_ (.CLK(clknet_leaf_38_clk),
    .D(_01168_),
    .Q(\dpath.alu.adder.in1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14957_ (.CLK(clknet_leaf_70_clk),
    .D(_01169_),
    .Q(\dpath.alu.adder.in1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_146_clk),
    .D(_01170_),
    .Q(\dpath.alu.adder.in1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14959_ (.CLK(clknet_leaf_70_clk),
    .D(_01171_),
    .Q(\dpath.alu.adder.in1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.CLK(clknet_leaf_70_clk),
    .D(_01172_),
    .Q(\dpath.alu.adder.in1[19] ));
 sky130_fd_sc_hd__dfxtp_4 _14961_ (.CLK(clknet_leaf_70_clk),
    .D(_01173_),
    .Q(\dpath.alu.adder.in1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.CLK(clknet_leaf_70_clk),
    .D(_01174_),
    .Q(\dpath.alu.adder.in1[21] ));
 sky130_fd_sc_hd__dfxtp_4 _14963_ (.CLK(clknet_leaf_70_clk),
    .D(_01175_),
    .Q(\dpath.alu.adder.in1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _14964_ (.CLK(clknet_leaf_70_clk),
    .D(_01176_),
    .Q(\dpath.alu.adder.in1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.CLK(clknet_leaf_70_clk),
    .D(_01177_),
    .Q(\dpath.alu.adder.in1[24] ));
 sky130_fd_sc_hd__dfxtp_4 _14966_ (.CLK(clknet_leaf_70_clk),
    .D(_01178_),
    .Q(\dpath.alu.adder.in1[25] ));
 sky130_fd_sc_hd__dfxtp_4 _14967_ (.CLK(clknet_leaf_70_clk),
    .D(_01179_),
    .Q(\dpath.alu.adder.in1[26] ));
 sky130_fd_sc_hd__dfxtp_4 _14968_ (.CLK(clknet_leaf_71_clk),
    .D(_01180_),
    .Q(\dpath.alu.adder.in1[27] ));
 sky130_fd_sc_hd__dfxtp_4 _14969_ (.CLK(clknet_leaf_71_clk),
    .D(_01181_),
    .Q(\dpath.alu.adder.in1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _14970_ (.CLK(clknet_leaf_75_clk),
    .D(_01182_),
    .Q(\dpath.alu.adder.in1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _14971_ (.CLK(clknet_leaf_70_clk),
    .D(_01183_),
    .Q(\dpath.alu.adder.in1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _14972_ (.CLK(clknet_leaf_71_clk),
    .D(_01184_),
    .Q(\dpath.alu.adder.in1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_65_clk),
    .D(net959),
    .Q(\dpath.csrw_out0.d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_92_clk),
    .D(net1055),
    .Q(\dpath.csrw_out0.d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_94_clk),
    .D(net965),
    .Q(\dpath.csrw_out0.d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.CLK(clknet_leaf_99_clk),
    .D(net957),
    .Q(\dpath.csrw_out0.d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.CLK(clknet_leaf_99_clk),
    .D(net1011),
    .Q(\dpath.csrw_out0.d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_99_clk),
    .D(net941),
    .Q(\dpath.csrw_out0.d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.CLK(clknet_leaf_99_clk),
    .D(net947),
    .Q(\dpath.csrw_out0.d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.CLK(clknet_leaf_96_clk),
    .D(net951),
    .Q(\dpath.csrw_out0.d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.CLK(clknet_leaf_95_clk),
    .D(net917),
    .Q(\dpath.csrw_out0.d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.CLK(clknet_leaf_97_clk),
    .D(net927),
    .Q(\dpath.csrw_out0.d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.CLK(clknet_leaf_96_clk),
    .D(net977),
    .Q(\dpath.csrw_out0.d[10] ));
 sky130_fd_sc_hd__dfxtp_4 _14984_ (.CLK(clknet_leaf_98_clk),
    .D(net963),
    .Q(\dpath.csrw_out0.d[11] ));
 sky130_fd_sc_hd__dfxtp_4 _14985_ (.CLK(clknet_leaf_100_clk),
    .D(net1043),
    .Q(\dpath.csrw_out0.d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.CLK(clknet_leaf_100_clk),
    .D(net897),
    .Q(\dpath.csrw_out0.d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14987_ (.CLK(clknet_leaf_98_clk),
    .D(net967),
    .Q(\dpath.csrw_out0.d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.CLK(clknet_leaf_96_clk),
    .D(net969),
    .Q(\dpath.csrw_out0.d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.CLK(clknet_leaf_106_clk),
    .D(net921),
    .Q(\dpath.csrw_out0.d[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.CLK(clknet_leaf_96_clk),
    .D(net971),
    .Q(\dpath.csrw_out0.d[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_105_clk),
    .D(net979),
    .Q(\dpath.csrw_out0.d[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_97_clk),
    .D(net935),
    .Q(\dpath.csrw_out0.d[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.CLK(clknet_leaf_99_clk),
    .D(net1033),
    .Q(\dpath.csrw_out0.d[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_99_clk),
    .D(net989),
    .Q(\dpath.csrw_out0.d[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_96_clk),
    .D(net929),
    .Q(\dpath.csrw_out0.d[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_92_clk),
    .D(net1013),
    .Q(\dpath.csrw_out0.d[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_92_clk),
    .D(net1049),
    .Q(\dpath.csrw_out0.d[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_93_clk),
    .D(net983),
    .Q(\dpath.csrw_out0.d[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_93_clk),
    .D(net975),
    .Q(\dpath.csrw_out0.d[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_93_clk),
    .D(net943),
    .Q(\dpath.csrw_out0.d[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_91_clk),
    .D(net997),
    .Q(\dpath.csrw_out0.d[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_91_clk),
    .D(net1037),
    .Q(\dpath.csrw_out0.d[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_91_clk),
    .D(net1067),
    .Q(\dpath.csrw_out0.d[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_92_clk),
    .D(net1603),
    .Q(\dpath.csrw_out0.d[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_175_clk),
    .D(_01217_),
    .Q(\dpath.sd_DX.q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.CLK(clknet_leaf_175_clk),
    .D(_01218_),
    .Q(\dpath.sd_DX.q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_174_clk),
    .D(_01219_),
    .Q(\dpath.sd_DX.q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_175_clk),
    .D(_01220_),
    .Q(\dpath.sd_DX.q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_175_clk),
    .D(_01221_),
    .Q(\dpath.sd_DX.q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.CLK(clknet_leaf_174_clk),
    .D(_01222_),
    .Q(\dpath.sd_DX.q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_175_clk),
    .D(_01223_),
    .Q(\dpath.sd_DX.q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_174_clk),
    .D(_01224_),
    .Q(\dpath.sd_DX.q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_170_clk),
    .D(_01225_),
    .Q(\dpath.sd_DX.q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_leaf_174_clk),
    .D(_01226_),
    .Q(\dpath.sd_DX.q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_154_clk),
    .D(_01227_),
    .Q(\dpath.sd_DX.q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_170_clk),
    .D(_01228_),
    .Q(\dpath.sd_DX.q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.CLK(clknet_leaf_170_clk),
    .D(_01229_),
    .Q(\dpath.sd_DX.q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.CLK(clknet_leaf_170_clk),
    .D(_01230_),
    .Q(\dpath.sd_DX.q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15019_ (.CLK(clknet_leaf_169_clk),
    .D(_01231_),
    .Q(\dpath.sd_DX.q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15020_ (.CLK(clknet_leaf_169_clk),
    .D(_01232_),
    .Q(\dpath.sd_DX.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15021_ (.CLK(clknet_leaf_120_clk),
    .D(_01233_),
    .Q(\dpath.sd_DX.q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.CLK(clknet_leaf_121_clk),
    .D(_01234_),
    .Q(\dpath.sd_DX.q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15023_ (.CLK(clknet_leaf_120_clk),
    .D(_01235_),
    .Q(\dpath.sd_DX.q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15024_ (.CLK(clknet_leaf_120_clk),
    .D(_01236_),
    .Q(\dpath.sd_DX.q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15025_ (.CLK(clknet_leaf_120_clk),
    .D(_01237_),
    .Q(\dpath.sd_DX.q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.CLK(clknet_leaf_120_clk),
    .D(_01238_),
    .Q(\dpath.sd_DX.q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15027_ (.CLK(clknet_leaf_120_clk),
    .D(_01239_),
    .Q(\dpath.sd_DX.q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15028_ (.CLK(clknet_leaf_119_clk),
    .D(_01240_),
    .Q(\dpath.sd_DX.q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15029_ (.CLK(clknet_leaf_119_clk),
    .D(_01241_),
    .Q(\dpath.sd_DX.q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15030_ (.CLK(clknet_leaf_119_clk),
    .D(_01242_),
    .Q(\dpath.sd_DX.q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15031_ (.CLK(clknet_leaf_140_clk),
    .D(_01243_),
    .Q(\dpath.sd_DX.q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15032_ (.CLK(clknet_leaf_136_clk),
    .D(_01244_),
    .Q(\dpath.sd_DX.q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.CLK(clknet_leaf_136_clk),
    .D(_01245_),
    .Q(\dpath.sd_DX.q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15034_ (.CLK(clknet_leaf_73_clk),
    .D(_01246_),
    .Q(\dpath.sd_DX.q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.CLK(clknet_leaf_143_clk),
    .D(_01247_),
    .Q(\dpath.sd_DX.q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.CLK(clknet_leaf_73_clk),
    .D(_01248_),
    .Q(\dpath.sd_DX.q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.CLK(clknet_leaf_23_clk),
    .D(_01249_),
    .Q(\dpath.RF.wdata[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15038_ (.CLK(clknet_leaf_23_clk),
    .D(_01250_),
    .Q(\dpath.RF.wdata[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15039_ (.CLK(clknet_leaf_26_clk),
    .D(_01251_),
    .Q(\dpath.RF.wdata[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15040_ (.CLK(clknet_leaf_184_clk),
    .D(_01252_),
    .Q(\dpath.RF.wdata[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15041_ (.CLK(clknet_leaf_180_clk),
    .D(_01253_),
    .Q(\dpath.RF.wdata[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15042_ (.CLK(clknet_leaf_178_clk),
    .D(_01254_),
    .Q(\dpath.RF.wdata[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15043_ (.CLK(clknet_leaf_2_clk),
    .D(_01255_),
    .Q(\dpath.RF.wdata[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.CLK(clknet_leaf_175_clk),
    .D(_01256_),
    .Q(\dpath.RF.wdata[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15045_ (.CLK(clknet_leaf_27_clk),
    .D(_01257_),
    .Q(\dpath.RF.wdata[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15046_ (.CLK(clknet_leaf_155_clk),
    .D(_01258_),
    .Q(\dpath.RF.wdata[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15047_ (.CLK(clknet_leaf_149_clk),
    .D(_01259_),
    .Q(\dpath.RF.wdata[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15048_ (.CLK(clknet_leaf_173_clk),
    .D(_01260_),
    .Q(\dpath.RF.wdata[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15049_ (.CLK(clknet_leaf_160_clk),
    .D(_01261_),
    .Q(\dpath.RF.wdata[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15050_ (.CLK(clknet_leaf_170_clk),
    .D(_01262_),
    .Q(\dpath.RF.wdata[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15051_ (.CLK(clknet_leaf_152_clk),
    .D(_01263_),
    .Q(\dpath.RF.wdata[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15052_ (.CLK(clknet_leaf_168_clk),
    .D(_01264_),
    .Q(\dpath.RF.wdata[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15053_ (.CLK(clknet_leaf_121_clk),
    .D(_01265_),
    .Q(\dpath.RF.wdata[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15054_ (.CLK(clknet_leaf_121_clk),
    .D(_01266_),
    .Q(\dpath.RF.wdata[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15055_ (.CLK(clknet_leaf_117_clk),
    .D(_01267_),
    .Q(\dpath.RF.wdata[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15056_ (.CLK(clknet_leaf_125_clk),
    .D(_01268_),
    .Q(\dpath.RF.wdata[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15057_ (.CLK(clknet_leaf_119_clk),
    .D(_01269_),
    .Q(\dpath.RF.wdata[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15058_ (.CLK(clknet_leaf_124_clk),
    .D(_01270_),
    .Q(\dpath.RF.wdata[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15059_ (.CLK(clknet_leaf_138_clk),
    .D(_01271_),
    .Q(\dpath.RF.wdata[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15060_ (.CLK(clknet_leaf_129_clk),
    .D(_01272_),
    .Q(\dpath.RF.wdata[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15061_ (.CLK(clknet_leaf_129_clk),
    .D(_01273_),
    .Q(\dpath.RF.wdata[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15062_ (.CLK(clknet_leaf_137_clk),
    .D(_01274_),
    .Q(\dpath.RF.wdata[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15063_ (.CLK(clknet_leaf_140_clk),
    .D(_01275_),
    .Q(\dpath.RF.wdata[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15064_ (.CLK(clknet_leaf_136_clk),
    .D(_01276_),
    .Q(\dpath.RF.wdata[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15065_ (.CLK(clknet_leaf_136_clk),
    .D(_01277_),
    .Q(\dpath.RF.wdata[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15066_ (.CLK(clknet_leaf_72_clk),
    .D(_01278_),
    .Q(\dpath.RF.wdata[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15067_ (.CLK(clknet_leaf_141_clk),
    .D(_01279_),
    .Q(\dpath.RF.wdata[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15068_ (.CLK(clknet_leaf_72_clk),
    .D(_01280_),
    .Q(\dpath.RF.wdata[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15069_ (.CLK(clknet_leaf_22_clk),
    .D(net1935),
    .Q(\dpath.RF.R[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15070_ (.CLK(clknet_leaf_24_clk),
    .D(net3123),
    .Q(\dpath.RF.R[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15071_ (.CLK(clknet_leaf_26_clk),
    .D(net3007),
    .Q(\dpath.RF.R[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15072_ (.CLK(clknet_leaf_187_clk),
    .D(net1831),
    .Q(\dpath.RF.R[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15073_ (.CLK(clknet_leaf_0_clk),
    .D(net1993),
    .Q(\dpath.RF.R[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15074_ (.CLK(clknet_leaf_158_clk),
    .D(net2369),
    .Q(\dpath.RF.R[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.CLK(clknet_leaf_4_clk),
    .D(net1917),
    .Q(\dpath.RF.R[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.CLK(clknet_leaf_185_clk),
    .D(net2949),
    .Q(\dpath.RF.R[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15077_ (.CLK(clknet_leaf_34_clk),
    .D(net1423),
    .Q(\dpath.RF.R[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15078_ (.CLK(clknet_leaf_155_clk),
    .D(net1785),
    .Q(\dpath.RF.R[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15079_ (.CLK(clknet_leaf_149_clk),
    .D(net1927),
    .Q(\dpath.RF.R[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15080_ (.CLK(clknet_leaf_176_clk),
    .D(net1877),
    .Q(\dpath.RF.R[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15081_ (.CLK(clknet_leaf_160_clk),
    .D(net2993),
    .Q(\dpath.RF.R[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15082_ (.CLK(clknet_leaf_171_clk),
    .D(net1823),
    .Q(\dpath.RF.R[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15083_ (.CLK(clknet_leaf_162_clk),
    .D(net2437),
    .Q(\dpath.RF.R[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15084_ (.CLK(clknet_leaf_168_clk),
    .D(net2155),
    .Q(\dpath.RF.R[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15085_ (.CLK(clknet_leaf_118_clk),
    .D(net1839),
    .Q(\dpath.RF.R[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.CLK(clknet_leaf_122_clk),
    .D(net1243),
    .Q(\dpath.RF.R[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.CLK(clknet_leaf_117_clk),
    .D(net1585),
    .Q(\dpath.RF.R[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.CLK(clknet_leaf_129_clk),
    .D(net1913),
    .Q(\dpath.RF.R[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.CLK(clknet_leaf_115_clk),
    .D(net1203),
    .Q(\dpath.RF.R[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.CLK(clknet_leaf_110_clk),
    .D(net2067),
    .Q(\dpath.RF.R[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.CLK(clknet_leaf_152_clk),
    .D(net1733),
    .Q(\dpath.RF.R[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.CLK(clknet_leaf_131_clk),
    .D(net2653),
    .Q(\dpath.RF.R[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.CLK(clknet_leaf_111_clk),
    .D(net1637),
    .Q(\dpath.RF.R[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.CLK(clknet_leaf_83_clk),
    .D(net1289),
    .Q(\dpath.RF.R[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15095_ (.CLK(clknet_leaf_141_clk),
    .D(net1419),
    .Q(\dpath.RF.R[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15096_ (.CLK(clknet_leaf_84_clk),
    .D(net1449),
    .Q(\dpath.RF.R[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15097_ (.CLK(clknet_leaf_73_clk),
    .D(net1307),
    .Q(\dpath.RF.R[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15098_ (.CLK(clknet_leaf_87_clk),
    .D(net1649),
    .Q(\dpath.RF.R[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15099_ (.CLK(clknet_leaf_143_clk),
    .D(net1347),
    .Q(\dpath.RF.R[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15100_ (.CLK(clknet_leaf_88_clk),
    .D(net1431),
    .Q(\dpath.RF.R[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15101_ (.CLK(clknet_leaf_57_clk),
    .D(_01313_),
    .Q(\dpath.csrr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.CLK(clknet_leaf_57_clk),
    .D(_01314_),
    .Q(\dpath.csrr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.CLK(clknet_leaf_57_clk),
    .D(_01315_),
    .Q(\dpath.csrr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.CLK(clknet_leaf_57_clk),
    .D(_01316_),
    .Q(\dpath.csrr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.CLK(clknet_leaf_57_clk),
    .D(_01317_),
    .Q(\dpath.csrr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.CLK(clknet_leaf_57_clk),
    .D(_01318_),
    .Q(\dpath.csrr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.CLK(clknet_leaf_57_clk),
    .D(_01319_),
    .Q(\dpath.csrr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.CLK(clknet_leaf_57_clk),
    .D(_01320_),
    .Q(\dpath.csrr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.CLK(clknet_leaf_57_clk),
    .D(_01321_),
    .Q(\dpath.csrr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.CLK(clknet_leaf_57_clk),
    .D(_01322_),
    .Q(\dpath.csrr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.CLK(clknet_leaf_57_clk),
    .D(_01323_),
    .Q(\dpath.csrr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.CLK(clknet_leaf_57_clk),
    .D(_01324_),
    .Q(\dpath.csrr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.CLK(clknet_leaf_57_clk),
    .D(_01325_),
    .Q(\dpath.csrr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.CLK(clknet_leaf_57_clk),
    .D(_01326_),
    .Q(\dpath.csrr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.CLK(clknet_leaf_57_clk),
    .D(_01327_),
    .Q(\dpath.csrr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.CLK(clknet_leaf_57_clk),
    .D(_01328_),
    .Q(\dpath.csrr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.CLK(clknet_leaf_58_clk),
    .D(_01329_),
    .Q(\dpath.csrr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.CLK(clknet_leaf_58_clk),
    .D(_01330_),
    .Q(\dpath.csrr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.CLK(clknet_leaf_58_clk),
    .D(_01331_),
    .Q(\dpath.csrr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.CLK(clknet_leaf_58_clk),
    .D(_01332_),
    .Q(\dpath.csrr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.CLK(clknet_leaf_58_clk),
    .D(_01333_),
    .Q(\dpath.csrr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15122_ (.CLK(clknet_leaf_59_clk),
    .D(_01334_),
    .Q(\dpath.csrr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15123_ (.CLK(clknet_leaf_59_clk),
    .D(_01335_),
    .Q(\dpath.csrr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15124_ (.CLK(clknet_leaf_59_clk),
    .D(_01336_),
    .Q(\dpath.csrr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15125_ (.CLK(clknet_leaf_58_clk),
    .D(_01337_),
    .Q(\dpath.csrr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15126_ (.CLK(clknet_leaf_59_clk),
    .D(_01338_),
    .Q(\dpath.csrr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15127_ (.CLK(clknet_leaf_58_clk),
    .D(_01339_),
    .Q(\dpath.csrr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15128_ (.CLK(clknet_leaf_59_clk),
    .D(_01340_),
    .Q(\dpath.csrr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15129_ (.CLK(clknet_leaf_59_clk),
    .D(_01341_),
    .Q(\dpath.csrr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15130_ (.CLK(clknet_leaf_59_clk),
    .D(_01342_),
    .Q(\dpath.csrr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15131_ (.CLK(clknet_leaf_59_clk),
    .D(_01343_),
    .Q(\dpath.csrr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15132_ (.CLK(clknet_leaf_59_clk),
    .D(_01344_),
    .Q(\dpath.csrr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15133_ (.CLK(clknet_leaf_13_clk),
    .D(_01345_),
    .Q(\dpath.btarg_DX.q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15134_ (.CLK(clknet_leaf_13_clk),
    .D(_01346_),
    .Q(\dpath.btarg_DX.q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15135_ (.CLK(clknet_leaf_15_clk),
    .D(_01347_),
    .Q(\dpath.btarg_DX.q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15136_ (.CLK(clknet_leaf_9_clk),
    .D(_01348_),
    .Q(\dpath.btarg_DX.q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15137_ (.CLK(clknet_leaf_5_clk),
    .D(_01349_),
    .Q(\dpath.btarg_DX.q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15138_ (.CLK(clknet_leaf_4_clk),
    .D(_01350_),
    .Q(\dpath.btarg_DX.q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15139_ (.CLK(clknet_leaf_4_clk),
    .D(_01351_),
    .Q(\dpath.btarg_DX.q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15140_ (.CLK(clknet_leaf_6_clk),
    .D(_01352_),
    .Q(\dpath.btarg_DX.q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15141_ (.CLK(clknet_leaf_9_clk),
    .D(_01353_),
    .Q(\dpath.btarg_DX.q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15142_ (.CLK(clknet_leaf_5_clk),
    .D(_01354_),
    .Q(\dpath.btarg_DX.q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15143_ (.CLK(clknet_leaf_9_clk),
    .D(_01355_),
    .Q(\dpath.btarg_DX.q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15144_ (.CLK(clknet_leaf_6_clk),
    .D(_01356_),
    .Q(\dpath.btarg_DX.q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15145_ (.CLK(clknet_leaf_7_clk),
    .D(_01357_),
    .Q(\dpath.btarg_DX.q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15146_ (.CLK(clknet_leaf_7_clk),
    .D(_01358_),
    .Q(\dpath.btarg_DX.q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15147_ (.CLK(clknet_leaf_7_clk),
    .D(_01359_),
    .Q(\dpath.btarg_DX.q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15148_ (.CLK(clknet_leaf_7_clk),
    .D(_01360_),
    .Q(\dpath.btarg_DX.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15149_ (.CLK(clknet_leaf_8_clk),
    .D(_01361_),
    .Q(\dpath.btarg_DX.q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15150_ (.CLK(clknet_leaf_8_clk),
    .D(_01362_),
    .Q(\dpath.btarg_DX.q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15151_ (.CLK(clknet_leaf_9_clk),
    .D(_01363_),
    .Q(\dpath.btarg_DX.q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15152_ (.CLK(clknet_leaf_9_clk),
    .D(_01364_),
    .Q(\dpath.btarg_DX.q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15153_ (.CLK(clknet_leaf_11_clk),
    .D(_01365_),
    .Q(\dpath.btarg_DX.q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15154_ (.CLK(clknet_leaf_11_clk),
    .D(_01366_),
    .Q(\dpath.btarg_DX.q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15155_ (.CLK(clknet_leaf_11_clk),
    .D(_01367_),
    .Q(\dpath.btarg_DX.q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15156_ (.CLK(clknet_leaf_12_clk),
    .D(_01368_),
    .Q(\dpath.btarg_DX.q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15157_ (.CLK(clknet_leaf_12_clk),
    .D(_01369_),
    .Q(\dpath.btarg_DX.q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15158_ (.CLK(clknet_leaf_13_clk),
    .D(_01370_),
    .Q(\dpath.btarg_DX.q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15159_ (.CLK(clknet_leaf_15_clk),
    .D(_01371_),
    .Q(\dpath.btarg_DX.q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15160_ (.CLK(clknet_leaf_14_clk),
    .D(_01372_),
    .Q(\dpath.btarg_DX.q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15161_ (.CLK(clknet_leaf_16_clk),
    .D(_01373_),
    .Q(\dpath.btarg_DX.q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15162_ (.CLK(clknet_leaf_16_clk),
    .D(_01374_),
    .Q(\dpath.btarg_DX.q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15163_ (.CLK(clknet_leaf_17_clk),
    .D(_01375_),
    .Q(\dpath.btarg_DX.q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15164_ (.CLK(clknet_leaf_14_clk),
    .D(_01376_),
    .Q(\dpath.btarg_DX.q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15165_ (.CLK(clknet_leaf_185_clk),
    .D(_01377_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_2 _15166_ (.CLK(clknet_leaf_185_clk),
    .D(_01378_),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_2 _15167_ (.CLK(clknet_leaf_185_clk),
    .D(_01379_),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _15168_ (.CLK(clknet_leaf_185_clk),
    .D(_01380_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_1 _15169_ (.CLK(clknet_leaf_185_clk),
    .D(_01381_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_2 _15170_ (.CLK(clknet_leaf_175_clk),
    .D(_01382_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_1 _15171_ (.CLK(clknet_leaf_185_clk),
    .D(_01383_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_2 _15172_ (.CLK(clknet_leaf_175_clk),
    .D(_01384_),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_2 _15173_ (.CLK(clknet_leaf_174_clk),
    .D(_01385_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_2 _15174_ (.CLK(clknet_leaf_174_clk),
    .D(_01386_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_2 _15175_ (.CLK(clknet_leaf_174_clk),
    .D(_01387_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _15176_ (.CLK(clknet_leaf_174_clk),
    .D(_01388_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_2 _15177_ (.CLK(clknet_leaf_174_clk),
    .D(_01389_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_2 _15178_ (.CLK(clknet_leaf_171_clk),
    .D(_01390_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_2 _15179_ (.CLK(clknet_leaf_170_clk),
    .D(_01391_),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_2 _15180_ (.CLK(clknet_leaf_169_clk),
    .D(_01392_),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_2 _15181_ (.CLK(clknet_leaf_120_clk),
    .D(_01393_),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_2 _15182_ (.CLK(clknet_leaf_169_clk),
    .D(_01394_),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_2 _15183_ (.CLK(clknet_leaf_119_clk),
    .D(_01395_),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_2 _15184_ (.CLK(clknet_leaf_169_clk),
    .D(_01396_),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_2 _15185_ (.CLK(clknet_leaf_119_clk),
    .D(_01397_),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_2 _15186_ (.CLK(clknet_leaf_119_clk),
    .D(_01398_),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_2 _15187_ (.CLK(clknet_leaf_121_clk),
    .D(_01399_),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_2 _15188_ (.CLK(clknet_leaf_120_clk),
    .D(_01400_),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_2 _15189_ (.CLK(clknet_leaf_119_clk),
    .D(_01401_),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_2 _15190_ (.CLK(clknet_leaf_119_clk),
    .D(_01402_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_2 _15191_ (.CLK(clknet_leaf_151_clk),
    .D(_01403_),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_4 _15192_ (.CLK(clknet_leaf_136_clk),
    .D(_01404_),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_4 _15193_ (.CLK(clknet_leaf_136_clk),
    .D(_01405_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_4 _15194_ (.CLK(clknet_leaf_73_clk),
    .D(_01406_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_2 _15195_ (.CLK(clknet_leaf_141_clk),
    .D(_01407_),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_4 _15196_ (.CLK(clknet_leaf_136_clk),
    .D(_01408_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_4 _15197_ (.CLK(clknet_leaf_49_clk),
    .D(_01409_),
    .Q(\dpath.alu.adder.in0[0] ));
 sky130_fd_sc_hd__dfxtp_4 _15198_ (.CLK(clknet_leaf_45_clk),
    .D(_01410_),
    .Q(\dpath.alu.adder.in0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15199_ (.CLK(clknet_leaf_45_clk),
    .D(_01411_),
    .Q(\dpath.alu.adder.in0[2] ));
 sky130_fd_sc_hd__dfxtp_4 _15200_ (.CLK(clknet_leaf_18_clk),
    .D(_01412_),
    .Q(\dpath.alu.adder.in0[3] ));
 sky130_fd_sc_hd__dfxtp_4 _15201_ (.CLK(clknet_leaf_18_clk),
    .D(_01413_),
    .Q(\dpath.alu.adder.in0[4] ));
 sky130_fd_sc_hd__dfxtp_4 _15202_ (.CLK(clknet_leaf_18_clk),
    .D(net1339),
    .Q(\dpath.alu.adder.in0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15203_ (.CLK(clknet_leaf_18_clk),
    .D(_01415_),
    .Q(\dpath.alu.adder.in0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15204_ (.CLK(clknet_leaf_18_clk),
    .D(_01416_),
    .Q(\dpath.alu.adder.in0[7] ));
 sky130_fd_sc_hd__dfxtp_4 _15205_ (.CLK(clknet_leaf_18_clk),
    .D(_01417_),
    .Q(\dpath.alu.adder.in0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15206_ (.CLK(clknet_leaf_19_clk),
    .D(net3229),
    .Q(\dpath.alu.adder.in0[9] ));
 sky130_fd_sc_hd__dfxtp_4 _15207_ (.CLK(clknet_leaf_19_clk),
    .D(_01419_),
    .Q(\dpath.alu.adder.in0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15208_ (.CLK(clknet_leaf_19_clk),
    .D(net3359),
    .Q(\dpath.alu.adder.in0[11] ));
 sky130_fd_sc_hd__dfxtp_4 _15209_ (.CLK(clknet_leaf_19_clk),
    .D(_01421_),
    .Q(\dpath.alu.adder.in0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15210_ (.CLK(clknet_leaf_19_clk),
    .D(_01422_),
    .Q(\dpath.alu.adder.in0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15211_ (.CLK(clknet_leaf_30_clk),
    .D(_01423_),
    .Q(\dpath.alu.adder.in0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15212_ (.CLK(clknet_leaf_30_clk),
    .D(_01424_),
    .Q(\dpath.alu.adder.in0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15213_ (.CLK(clknet_leaf_23_clk),
    .D(_01425_),
    .Q(\dpath.alu.adder.in0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15214_ (.CLK(clknet_leaf_44_clk),
    .D(_01426_),
    .Q(\dpath.alu.adder.in0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15215_ (.CLK(clknet_leaf_40_clk),
    .D(_01427_),
    .Q(\dpath.alu.adder.in0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15216_ (.CLK(clknet_leaf_40_clk),
    .D(_01428_),
    .Q(\dpath.alu.adder.in0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15217_ (.CLK(clknet_leaf_40_clk),
    .D(_01429_),
    .Q(\dpath.alu.adder.in0[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15218_ (.CLK(clknet_leaf_40_clk),
    .D(_01430_),
    .Q(\dpath.alu.adder.in0[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15219_ (.CLK(clknet_leaf_40_clk),
    .D(_01431_),
    .Q(\dpath.alu.adder.in0[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15220_ (.CLK(clknet_leaf_40_clk),
    .D(_01432_),
    .Q(\dpath.alu.adder.in0[23] ));
 sky130_fd_sc_hd__dfxtp_4 _15221_ (.CLK(clknet_leaf_41_clk),
    .D(_01433_),
    .Q(\dpath.alu.adder.in0[24] ));
 sky130_fd_sc_hd__dfxtp_4 _15222_ (.CLK(clknet_leaf_40_clk),
    .D(_01434_),
    .Q(\dpath.alu.adder.in0[25] ));
 sky130_fd_sc_hd__dfxtp_4 _15223_ (.CLK(clknet_leaf_19_clk),
    .D(_01435_),
    .Q(\dpath.alu.adder.in0[26] ));
 sky130_fd_sc_hd__dfxtp_4 _15224_ (.CLK(clknet_leaf_19_clk),
    .D(net3340),
    .Q(\dpath.alu.adder.in0[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15225_ (.CLK(clknet_leaf_41_clk),
    .D(_01437_),
    .Q(\dpath.alu.adder.in0[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15226_ (.CLK(clknet_leaf_19_clk),
    .D(net3440),
    .Q(\dpath.alu.adder.in0[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15227_ (.CLK(clknet_leaf_18_clk),
    .D(net3338),
    .Q(\dpath.alu.adder.in0[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15228_ (.CLK(clknet_leaf_18_clk),
    .D(net3185),
    .Q(\dpath.alu.adder.in0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15229_ (.CLK(clknet_leaf_66_clk),
    .D(net1141),
    .Q(\dpath.csrw_out_MW.d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15230_ (.CLK(clknet_leaf_91_clk),
    .D(net2621),
    .Q(\dpath.csrw_out_MW.d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15231_ (.CLK(clknet_leaf_95_clk),
    .D(net3171),
    .Q(\dpath.csrw_out_MW.d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15232_ (.CLK(clknet_leaf_100_clk),
    .D(net3195),
    .Q(\dpath.csrw_out_MW.d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15233_ (.CLK(clknet_leaf_99_clk),
    .D(_01445_),
    .Q(\dpath.csrw_out_MW.d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15234_ (.CLK(clknet_leaf_100_clk),
    .D(net2093),
    .Q(\dpath.csrw_out_MW.d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15235_ (.CLK(clknet_leaf_100_clk),
    .D(_01447_),
    .Q(\dpath.csrw_out_MW.d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15236_ (.CLK(clknet_leaf_95_clk),
    .D(net3179),
    .Q(\dpath.csrw_out_MW.d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15237_ (.CLK(clknet_leaf_86_clk),
    .D(net903),
    .Q(\dpath.csrw_out_MW.d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15238_ (.CLK(clknet_leaf_96_clk),
    .D(_01450_),
    .Q(\dpath.csrw_out_MW.d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15239_ (.CLK(clknet_leaf_101_clk),
    .D(net1019),
    .Q(\dpath.csrw_out_MW.d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15240_ (.CLK(clknet_leaf_100_clk),
    .D(net1971),
    .Q(\dpath.csrw_out_MW.d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15241_ (.CLK(clknet_leaf_100_clk),
    .D(net899),
    .Q(\dpath.csrw_out_MW.d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15242_ (.CLK(clknet_leaf_102_clk),
    .D(net1003),
    .Q(\dpath.csrw_out_MW.d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15243_ (.CLK(clknet_leaf_100_clk),
    .D(net993),
    .Q(\dpath.csrw_out_MW.d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15244_ (.CLK(clknet_leaf_101_clk),
    .D(net981),
    .Q(\dpath.csrw_out_MW.d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15245_ (.CLK(clknet_leaf_105_clk),
    .D(net1017),
    .Q(\dpath.csrw_out_MW.d[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15246_ (.CLK(clknet_leaf_86_clk),
    .D(net905),
    .Q(\dpath.csrw_out_MW.d[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15247_ (.CLK(clknet_leaf_105_clk),
    .D(net985),
    .Q(\dpath.csrw_out_MW.d[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15248_ (.CLK(clknet_leaf_96_clk),
    .D(net931),
    .Q(\dpath.csrw_out_MW.d[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15249_ (.CLK(clknet_leaf_99_clk),
    .D(net955),
    .Q(\dpath.csrw_out_MW.d[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15250_ (.CLK(clknet_leaf_99_clk),
    .D(net949),
    .Q(\dpath.csrw_out_MW.d[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15251_ (.CLK(clknet_leaf_95_clk),
    .D(net953),
    .Q(\dpath.csrw_out_MW.d[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15252_ (.CLK(clknet_leaf_91_clk),
    .D(net1029),
    .Q(\dpath.csrw_out_MW.d[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15253_ (.CLK(clknet_leaf_91_clk),
    .D(net937),
    .Q(\dpath.csrw_out_MW.d[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15254_ (.CLK(clknet_leaf_93_clk),
    .D(net919),
    .Q(\dpath.csrw_out_MW.d[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15255_ (.CLK(clknet_leaf_90_clk),
    .D(net995),
    .Q(\dpath.csrw_out_MW.d[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15256_ (.CLK(clknet_leaf_90_clk),
    .D(net1005),
    .Q(\dpath.csrw_out_MW.d[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15257_ (.CLK(clknet_leaf_91_clk),
    .D(net939),
    .Q(\dpath.csrw_out_MW.d[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15258_ (.CLK(clknet_leaf_91_clk),
    .D(net3063),
    .Q(\dpath.csrw_out_MW.d[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15259_ (.CLK(clknet_leaf_89_clk),
    .D(net1009),
    .Q(\dpath.csrw_out_MW.d[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15260_ (.CLK(clknet_leaf_89_clk),
    .D(net901),
    .Q(\dpath.csrw_out_MW.d[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15261_ (.CLK(clknet_leaf_22_clk),
    .D(net3057),
    .Q(\dpath.RF.R[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15262_ (.CLK(clknet_leaf_3_clk),
    .D(net2251),
    .Q(\dpath.RF.R[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15263_ (.CLK(clknet_leaf_29_clk),
    .D(net1939),
    .Q(\dpath.RF.R[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15264_ (.CLK(clknet_leaf_186_clk),
    .D(net3157),
    .Q(\dpath.RF.R[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15265_ (.CLK(clknet_leaf_0_clk),
    .D(net2907),
    .Q(\dpath.RF.R[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15266_ (.CLK(clknet_leaf_158_clk),
    .D(net3017),
    .Q(\dpath.RF.R[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15267_ (.CLK(clknet_leaf_3_clk),
    .D(net2781),
    .Q(\dpath.RF.R[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15268_ (.CLK(clknet_leaf_175_clk),
    .D(net2833),
    .Q(\dpath.RF.R[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15269_ (.CLK(clknet_leaf_35_clk),
    .D(net2313),
    .Q(\dpath.RF.R[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15270_ (.CLK(clknet_leaf_155_clk),
    .D(net2923),
    .Q(\dpath.RF.R[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15271_ (.CLK(clknet_leaf_148_clk),
    .D(net3045),
    .Q(\dpath.RF.R[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15272_ (.CLK(clknet_leaf_173_clk),
    .D(net1601),
    .Q(\dpath.RF.R[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15273_ (.CLK(clknet_leaf_160_clk),
    .D(net2741),
    .Q(\dpath.RF.R[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15274_ (.CLK(clknet_leaf_171_clk),
    .D(net3191),
    .Q(\dpath.RF.R[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15275_ (.CLK(clknet_leaf_152_clk),
    .D(net2179),
    .Q(\dpath.RF.R[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15276_ (.CLK(clknet_leaf_167_clk),
    .D(net1843),
    .Q(\dpath.RF.R[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15277_ (.CLK(clknet_leaf_118_clk),
    .D(net2209),
    .Q(\dpath.RF.R[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15278_ (.CLK(clknet_leaf_121_clk),
    .D(net2405),
    .Q(\dpath.RF.R[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15279_ (.CLK(clknet_leaf_116_clk),
    .D(net3065),
    .Q(\dpath.RF.R[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15280_ (.CLK(clknet_leaf_129_clk),
    .D(net2301),
    .Q(\dpath.RF.R[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15281_ (.CLK(clknet_leaf_108_clk),
    .D(net2507),
    .Q(\dpath.RF.R[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15282_ (.CLK(clknet_leaf_109_clk),
    .D(net2217),
    .Q(\dpath.RF.R[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15283_ (.CLK(clknet_leaf_152_clk),
    .D(net1847),
    .Q(\dpath.RF.R[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15284_ (.CLK(clknet_leaf_131_clk),
    .D(net2627),
    .Q(\dpath.RF.R[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15285_ (.CLK(clknet_leaf_103_clk),
    .D(net1521),
    .Q(\dpath.RF.R[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15286_ (.CLK(clknet_leaf_83_clk),
    .D(net2969),
    .Q(\dpath.RF.R[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15287_ (.CLK(clknet_leaf_144_clk),
    .D(net1345),
    .Q(\dpath.RF.R[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15288_ (.CLK(clknet_leaf_84_clk),
    .D(net2505),
    .Q(\dpath.RF.R[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15289_ (.CLK(clknet_leaf_73_clk),
    .D(net1859),
    .Q(\dpath.RF.R[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15290_ (.CLK(clknet_leaf_87_clk),
    .D(net2041),
    .Q(\dpath.RF.R[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15291_ (.CLK(clknet_leaf_143_clk),
    .D(net1573),
    .Q(\dpath.RF.R[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15292_ (.CLK(clknet_leaf_88_clk),
    .D(net1665),
    .Q(\dpath.RF.R[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15293_ (.CLK(clknet_leaf_43_clk),
    .D(_01505_),
    .Q(\ctrl.val_M ));
 sky130_fd_sc_hd__dfxtp_1 _15294_ (.CLK(clknet_leaf_49_clk),
    .D(_01506_),
    .Q(\dpath.inst_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15295_ (.CLK(clknet_leaf_49_clk),
    .D(net3234),
    .Q(\dpath.inst_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15296_ (.CLK(clknet_leaf_16_clk),
    .D(_01508_),
    .Q(\dpath.inst_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15297_ (.CLK(clknet_leaf_15_clk),
    .D(net3232),
    .Q(\dpath.inst_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15298_ (.CLK(clknet_leaf_5_clk),
    .D(net3239),
    .Q(\dpath.inst_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15299_ (.CLK(clknet_leaf_4_clk),
    .D(_01511_),
    .Q(\dpath.inst_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15300_ (.CLK(clknet_leaf_5_clk),
    .D(net3298),
    .Q(\dpath.inst_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15301_ (.CLK(clknet_leaf_5_clk),
    .D(net3278),
    .Q(\dpath.inst_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15302_ (.CLK(clknet_leaf_9_clk),
    .D(net3287),
    .Q(\dpath.inst_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15303_ (.CLK(clknet_leaf_6_clk),
    .D(_01515_),
    .Q(\dpath.inst_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15304_ (.CLK(clknet_leaf_9_clk),
    .D(net3275),
    .Q(\dpath.inst_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15305_ (.CLK(clknet_leaf_6_clk),
    .D(_01517_),
    .Q(\dpath.inst_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15306_ (.CLK(clknet_leaf_7_clk),
    .D(net3302),
    .Q(\dpath.inst_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15307_ (.CLK(clknet_leaf_7_clk),
    .D(net3296),
    .Q(\dpath.inst_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15308_ (.CLK(clknet_leaf_7_clk),
    .D(net3292),
    .Q(\dpath.inst_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15309_ (.CLK(clknet_leaf_7_clk),
    .D(net3242),
    .Q(\dpath.inst_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15310_ (.CLK(clknet_leaf_8_clk),
    .D(net3266),
    .Q(\dpath.inst_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15311_ (.CLK(clknet_leaf_8_clk),
    .D(net3222),
    .Q(\dpath.inst_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15312_ (.CLK(clknet_leaf_11_clk),
    .D(net3326),
    .Q(\dpath.inst_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15313_ (.CLK(clknet_leaf_8_clk),
    .D(net3324),
    .Q(\dpath.inst_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15314_ (.CLK(clknet_leaf_10_clk),
    .D(net3463),
    .Q(\dpath.inst_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15315_ (.CLK(clknet_leaf_10_clk),
    .D(net3456),
    .Q(\dpath.inst_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15316_ (.CLK(clknet_leaf_11_clk),
    .D(net3467),
    .Q(\dpath.inst_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15317_ (.CLK(clknet_leaf_12_clk),
    .D(net3469),
    .Q(\dpath.inst_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15318_ (.CLK(clknet_leaf_12_clk),
    .D(_01530_),
    .Q(\dpath.inst_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15319_ (.CLK(clknet_leaf_13_clk),
    .D(_01531_),
    .Q(\dpath.inst_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15320_ (.CLK(clknet_leaf_15_clk),
    .D(_01532_),
    .Q(\dpath.inst_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15321_ (.CLK(clknet_leaf_14_clk),
    .D(_01533_),
    .Q(\dpath.inst_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15322_ (.CLK(clknet_leaf_18_clk),
    .D(net3402),
    .Q(\dpath.inst_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15323_ (.CLK(clknet_leaf_18_clk),
    .D(_01535_),
    .Q(\dpath.inst_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15324_ (.CLK(clknet_leaf_18_clk),
    .D(net3284),
    .Q(\dpath.inst_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15325_ (.CLK(clknet_leaf_14_clk),
    .D(_01537_),
    .Q(\dpath.inst_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15326_ (.CLK(clknet_leaf_50_clk),
    .D(_01538_),
    .Q(\ctrl.d2c_inst[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15327_ (.CLK(clknet_leaf_50_clk),
    .D(_01539_),
    .Q(\ctrl.d2c_inst[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15328_ (.CLK(clknet_leaf_50_clk),
    .D(_01540_),
    .Q(\ctrl.d2c_inst[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15329_ (.CLK(clknet_leaf_50_clk),
    .D(_01541_),
    .Q(\ctrl.d2c_inst[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15330_ (.CLK(clknet_leaf_51_clk),
    .D(_01542_),
    .Q(\ctrl.d2c_inst[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15331_ (.CLK(clknet_leaf_50_clk),
    .D(_01543_),
    .Q(\ctrl.d2c_inst[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15332_ (.CLK(clknet_leaf_51_clk),
    .D(_01544_),
    .Q(\ctrl.d2c_inst[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15333_ (.CLK(clknet_leaf_51_clk),
    .D(_01545_),
    .Q(\ctrl.d2c_inst[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15334_ (.CLK(clknet_leaf_51_clk),
    .D(_01546_),
    .Q(\ctrl.d2c_inst[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15335_ (.CLK(clknet_leaf_55_clk),
    .D(_01547_),
    .Q(\ctrl.d2c_inst[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15336_ (.CLK(clknet_leaf_51_clk),
    .D(_01548_),
    .Q(\ctrl.d2c_inst[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15337_ (.CLK(clknet_leaf_51_clk),
    .D(_01549_),
    .Q(\ctrl.d2c_inst[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15338_ (.CLK(clknet_leaf_52_clk),
    .D(_01550_),
    .Q(\ctrl.d2c_inst[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15339_ (.CLK(clknet_leaf_52_clk),
    .D(_01551_),
    .Q(\ctrl.d2c_inst[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15340_ (.CLK(clknet_leaf_51_clk),
    .D(_01552_),
    .Q(\ctrl.d2c_inst[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15341_ (.CLK(clknet_leaf_50_clk),
    .D(_01553_),
    .Q(\ctrl.d2c_inst[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15342_ (.CLK(clknet_leaf_50_clk),
    .D(_01554_),
    .Q(\ctrl.d2c_inst[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15343_ (.CLK(clknet_leaf_49_clk),
    .D(_01555_),
    .Q(\ctrl.d2c_inst[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15344_ (.CLK(clknet_leaf_49_clk),
    .D(_01556_),
    .Q(\ctrl.d2c_inst[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15345_ (.CLK(clknet_leaf_50_clk),
    .D(_01557_),
    .Q(\ctrl.d2c_inst[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15346_ (.CLK(clknet_leaf_48_clk),
    .D(_01558_),
    .Q(\ctrl.d2c_inst[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15347_ (.CLK(clknet_leaf_49_clk),
    .D(_01559_),
    .Q(\ctrl.d2c_inst[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15348_ (.CLK(clknet_leaf_48_clk),
    .D(_01560_),
    .Q(\ctrl.d2c_inst[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15349_ (.CLK(clknet_leaf_46_clk),
    .D(_01561_),
    .Q(\ctrl.d2c_inst[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15350_ (.CLK(clknet_leaf_46_clk),
    .D(_01562_),
    .Q(\ctrl.d2c_inst[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15351_ (.CLK(clknet_leaf_53_clk),
    .D(_01563_),
    .Q(\ctrl.d2c_inst[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15352_ (.CLK(clknet_leaf_54_clk),
    .D(_01564_),
    .Q(\ctrl.d2c_inst[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15353_ (.CLK(clknet_leaf_55_clk),
    .D(_01565_),
    .Q(\ctrl.d2c_inst[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15354_ (.CLK(clknet_leaf_55_clk),
    .D(_01566_),
    .Q(\ctrl.d2c_inst[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15355_ (.CLK(clknet_leaf_54_clk),
    .D(_01567_),
    .Q(\ctrl.d2c_inst[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15356_ (.CLK(clknet_leaf_54_clk),
    .D(_01568_),
    .Q(\ctrl.d2c_inst[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15357_ (.CLK(clknet_leaf_52_clk),
    .D(_01569_),
    .Q(\ctrl.d2c_inst[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15358_ (.CLK(clknet_leaf_23_clk),
    .D(net1813),
    .Q(\dpath.RF.R[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.CLK(clknet_leaf_24_clk),
    .D(net1779),
    .Q(\dpath.RF.R[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15360_ (.CLK(clknet_leaf_26_clk),
    .D(net2071),
    .Q(\dpath.RF.R[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15361_ (.CLK(clknet_leaf_182_clk),
    .D(net2051),
    .Q(\dpath.RF.R[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15362_ (.CLK(clknet_leaf_181_clk),
    .D(net1845),
    .Q(\dpath.RF.R[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15363_ (.CLK(clknet_leaf_158_clk),
    .D(net1789),
    .Q(\dpath.RF.R[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15364_ (.CLK(clknet_leaf_3_clk),
    .D(net1919),
    .Q(\dpath.RF.R[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15365_ (.CLK(clknet_leaf_185_clk),
    .D(net1543),
    .Q(\dpath.RF.R[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15366_ (.CLK(clknet_leaf_35_clk),
    .D(net3027),
    .Q(\dpath.RF.R[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15367_ (.CLK(clknet_leaf_153_clk),
    .D(net1235),
    .Q(\dpath.RF.R[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15368_ (.CLK(clknet_leaf_148_clk),
    .D(net1909),
    .Q(\dpath.RF.R[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15369_ (.CLK(clknet_leaf_173_clk),
    .D(net1367),
    .Q(\dpath.RF.R[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.CLK(clknet_leaf_160_clk),
    .D(net2415),
    .Q(\dpath.RF.R[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.CLK(clknet_leaf_171_clk),
    .D(net1355),
    .Q(\dpath.RF.R[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.CLK(clknet_leaf_162_clk),
    .D(net1477),
    .Q(\dpath.RF.R[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.CLK(clknet_leaf_168_clk),
    .D(net1741),
    .Q(\dpath.RF.R[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.CLK(clknet_leaf_118_clk),
    .D(net1663),
    .Q(\dpath.RF.R[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15375_ (.CLK(clknet_leaf_122_clk),
    .D(net1269),
    .Q(\dpath.RF.R[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.CLK(clknet_leaf_116_clk),
    .D(net2763),
    .Q(\dpath.RF.R[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.CLK(clknet_leaf_129_clk),
    .D(net1591),
    .Q(\dpath.RF.R[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15378_ (.CLK(clknet_leaf_108_clk),
    .D(net1273),
    .Q(\dpath.RF.R[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15379_ (.CLK(clknet_leaf_109_clk),
    .D(net1343),
    .Q(\dpath.RF.R[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15380_ (.CLK(clknet_leaf_139_clk),
    .D(net1447),
    .Q(\dpath.RF.R[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15381_ (.CLK(clknet_leaf_131_clk),
    .D(net2911),
    .Q(\dpath.RF.R[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15382_ (.CLK(clknet_leaf_103_clk),
    .D(net1739),
    .Q(\dpath.RF.R[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15383_ (.CLK(clknet_leaf_83_clk),
    .D(net2223),
    .Q(\dpath.RF.R[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15384_ (.CLK(clknet_leaf_141_clk),
    .D(net1211),
    .Q(\dpath.RF.R[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15385_ (.CLK(clknet_leaf_84_clk),
    .D(net2261),
    .Q(\dpath.RF.R[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15386_ (.CLK(clknet_leaf_78_clk),
    .D(net2497),
    .Q(\dpath.RF.R[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15387_ (.CLK(clknet_leaf_87_clk),
    .D(net2227),
    .Q(\dpath.RF.R[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15388_ (.CLK(clknet_leaf_143_clk),
    .D(net1849),
    .Q(\dpath.RF.R[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15389_ (.CLK(clknet_leaf_89_clk),
    .D(net1263),
    .Q(\dpath.RF.R[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15390_ (.CLK(clknet_leaf_20_clk),
    .D(net2663),
    .Q(\dpath.RF.R[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15391_ (.CLK(clknet_leaf_156_clk),
    .D(net2171),
    .Q(\dpath.RF.R[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15392_ (.CLK(clknet_leaf_31_clk),
    .D(net2059),
    .Q(\dpath.RF.R[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15393_ (.CLK(clknet_leaf_180_clk),
    .D(net2229),
    .Q(\dpath.RF.R[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15394_ (.CLK(clknet_leaf_1_clk),
    .D(net2539),
    .Q(\dpath.RF.R[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15395_ (.CLK(clknet_leaf_157_clk),
    .D(net2425),
    .Q(\dpath.RF.R[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15396_ (.CLK(clknet_leaf_2_clk),
    .D(net1537),
    .Q(\dpath.RF.R[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15397_ (.CLK(clknet_leaf_181_clk),
    .D(net1415),
    .Q(\dpath.RF.R[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15398_ (.CLK(clknet_leaf_32_clk),
    .D(net2219),
    .Q(\dpath.RF.R[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15399_ (.CLK(clknet_leaf_154_clk),
    .D(net1607),
    .Q(\dpath.RF.R[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15400_ (.CLK(clknet_leaf_35_clk),
    .D(net1095),
    .Q(\dpath.RF.R[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15401_ (.CLK(clknet_leaf_177_clk),
    .D(net1673),
    .Q(\dpath.RF.R[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15402_ (.CLK(clknet_leaf_165_clk),
    .D(net1699),
    .Q(\dpath.RF.R[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15403_ (.CLK(clknet_leaf_160_clk),
    .D(net2739),
    .Q(\dpath.RF.R[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15404_ (.CLK(clknet_leaf_152_clk),
    .D(net1805),
    .Q(\dpath.RF.R[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15405_ (.CLK(clknet_leaf_165_clk),
    .D(net1505),
    .Q(\dpath.RF.R[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15406_ (.CLK(clknet_leaf_124_clk),
    .D(net1301),
    .Q(\dpath.RF.R[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15407_ (.CLK(clknet_leaf_126_clk),
    .D(net2117),
    .Q(\dpath.RF.R[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15408_ (.CLK(clknet_leaf_131_clk),
    .D(net2503),
    .Q(\dpath.RF.R[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15409_ (.CLK(clknet_leaf_127_clk),
    .D(net1775),
    .Q(\dpath.RF.R[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15410_ (.CLK(clknet_leaf_114_clk),
    .D(net2615),
    .Q(\dpath.RF.R[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15411_ (.CLK(clknet_leaf_113_clk),
    .D(net2709),
    .Q(\dpath.RF.R[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15412_ (.CLK(clknet_leaf_138_clk),
    .D(net3053),
    .Q(\dpath.RF.R[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15413_ (.CLK(clknet_leaf_134_clk),
    .D(net1575),
    .Q(\dpath.RF.R[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15414_ (.CLK(clknet_leaf_132_clk),
    .D(net2365),
    .Q(\dpath.RF.R[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15415_ (.CLK(clknet_leaf_133_clk),
    .D(net1315),
    .Q(\dpath.RF.R[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15416_ (.CLK(clknet_leaf_148_clk),
    .D(net1715),
    .Q(\dpath.RF.R[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15417_ (.CLK(clknet_leaf_81_clk),
    .D(net2555),
    .Q(\dpath.RF.R[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15418_ (.CLK(clknet_leaf_75_clk),
    .D(net1703),
    .Q(\dpath.RF.R[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15419_ (.CLK(clknet_leaf_76_clk),
    .D(net2661),
    .Q(\dpath.RF.R[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15420_ (.CLK(clknet_leaf_143_clk),
    .D(net1679),
    .Q(\dpath.RF.R[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15421_ (.CLK(clknet_leaf_78_clk),
    .D(net2151),
    .Q(\dpath.RF.R[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15422_ (.CLK(clknet_leaf_50_clk),
    .D(_01634_),
    .Q(_00005_));
 sky130_fd_sc_hd__dfxtp_4 _15423_ (.CLK(clknet_leaf_12_clk),
    .D(net3227),
    .Q(_00006_));
 sky130_fd_sc_hd__dfxtp_4 _15424_ (.CLK(clknet_leaf_49_clk),
    .D(_01636_),
    .Q(_00007_));
 sky130_fd_sc_hd__dfxtp_4 _15425_ (.CLK(clknet_leaf_46_clk),
    .D(_01637_),
    .Q(_00008_));
 sky130_fd_sc_hd__dfxtp_4 _15426_ (.CLK(clknet_leaf_17_clk),
    .D(_01638_),
    .Q(_00009_));
 sky130_fd_sc_hd__dfxtp_1 _15427_ (.CLK(clknet_leaf_23_clk),
    .D(net2557),
    .Q(\dpath.RF.R[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15428_ (.CLK(clknet_leaf_24_clk),
    .D(net2393),
    .Q(\dpath.RF.R[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15429_ (.CLK(clknet_leaf_30_clk),
    .D(net1531),
    .Q(\dpath.RF.R[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15430_ (.CLK(clknet_leaf_180_clk),
    .D(net2565),
    .Q(\dpath.RF.R[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15431_ (.CLK(clknet_leaf_2_clk),
    .D(net1707),
    .Q(\dpath.RF.R[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15432_ (.CLK(clknet_leaf_158_clk),
    .D(net1557),
    .Q(\dpath.RF.R[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15433_ (.CLK(clknet_leaf_2_clk),
    .D(net1943),
    .Q(\dpath.RF.R[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15434_ (.CLK(clknet_leaf_180_clk),
    .D(net2551),
    .Q(\dpath.RF.R[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15435_ (.CLK(clknet_leaf_33_clk),
    .D(net2439),
    .Q(\dpath.RF.R[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15436_ (.CLK(clknet_leaf_154_clk),
    .D(net2165),
    .Q(\dpath.RF.R[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15437_ (.CLK(clknet_leaf_36_clk),
    .D(net1661),
    .Q(\dpath.RF.R[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15438_ (.CLK(clknet_leaf_177_clk),
    .D(net2929),
    .Q(\dpath.RF.R[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15439_ (.CLK(clknet_leaf_163_clk),
    .D(net1851),
    .Q(\dpath.RF.R[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15440_ (.CLK(clknet_leaf_160_clk),
    .D(net2029),
    .Q(\dpath.RF.R[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15441_ (.CLK(clknet_leaf_152_clk),
    .D(net2291),
    .Q(\dpath.RF.R[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15442_ (.CLK(clknet_leaf_164_clk),
    .D(net1777),
    .Q(\dpath.RF.R[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15443_ (.CLK(clknet_leaf_124_clk),
    .D(net1291),
    .Q(\dpath.RF.R[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15444_ (.CLK(clknet_leaf_126_clk),
    .D(net1619),
    .Q(\dpath.RF.R[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15445_ (.CLK(clknet_leaf_130_clk),
    .D(net1323),
    .Q(\dpath.RF.R[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15446_ (.CLK(clknet_leaf_127_clk),
    .D(net1407),
    .Q(\dpath.RF.R[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15447_ (.CLK(clknet_leaf_112_clk),
    .D(net1811),
    .Q(\dpath.RF.R[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15448_ (.CLK(clknet_leaf_112_clk),
    .D(net2015),
    .Q(\dpath.RF.R[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15449_ (.CLK(clknet_leaf_138_clk),
    .D(net2843),
    .Q(\dpath.RF.R[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15450_ (.CLK(clknet_leaf_135_clk),
    .D(net1225),
    .Q(\dpath.RF.R[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15451_ (.CLK(clknet_leaf_132_clk),
    .D(net1251),
    .Q(\dpath.RF.R[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15452_ (.CLK(clknet_leaf_134_clk),
    .D(net1333),
    .Q(\dpath.RF.R[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15453_ (.CLK(clknet_leaf_145_clk),
    .D(net1729),
    .Q(\dpath.RF.R[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15454_ (.CLK(clknet_leaf_81_clk),
    .D(net1611),
    .Q(\dpath.RF.R[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15455_ (.CLK(clknet_leaf_74_clk),
    .D(net1471),
    .Q(\dpath.RF.R[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15456_ (.CLK(clknet_leaf_76_clk),
    .D(net1725),
    .Q(\dpath.RF.R[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15457_ (.CLK(clknet_leaf_143_clk),
    .D(net1295),
    .Q(\dpath.RF.R[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15458_ (.CLK(clknet_leaf_77_clk),
    .D(net1257),
    .Q(\dpath.RF.R[30][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15459_ (.CLK(clknet_leaf_13_clk),
    .D(net3262),
    .Q(net228));
 sky130_fd_sc_hd__dfxtp_2 _15460_ (.CLK(clknet_leaf_13_clk),
    .D(net3528),
    .Q(net239));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_4 fanout1 (.A(_06815_),
    .X(net3719));
 sky130_fd_sc_hd__buf_4 fanout2 (.A(_06815_),
    .X(net3720));
 sky130_fd_sc_hd__buf_4 fanout3 (.A(_06814_),
    .X(net3721));
 sky130_fd_sc_hd__buf_8 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_16 fanout358 (.A(_06063_),
    .X(net358));
 sky130_fd_sc_hd__buf_12 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_12 fanout360 (.A(_06059_),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_8 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_8 fanout362 (.A(_01957_),
    .X(net362));
 sky130_fd_sc_hd__buf_6 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_8 fanout364 (.A(_06043_),
    .X(net364));
 sky130_fd_sc_hd__buf_4 fanout365 (.A(_02119_),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_8 fanout366 (.A(_02119_),
    .X(net366));
 sky130_fd_sc_hd__buf_8 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__buf_8 fanout368 (.A(_02116_),
    .X(net368));
 sky130_fd_sc_hd__buf_8 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_16 fanout370 (.A(_02115_),
    .X(net370));
 sky130_fd_sc_hd__buf_8 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_8 fanout372 (.A(_02097_),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_8 fanout373 (.A(_02028_),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_4 fanout374 (.A(_02028_),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_16 fanout375 (.A(_01685_),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_16 fanout376 (.A(_01685_),
    .X(net376));
 sky130_fd_sc_hd__buf_6 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_16 fanout378 (.A(_06056_),
    .X(net378));
 sky130_fd_sc_hd__buf_8 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_16 fanout380 (.A(_06042_),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_16 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_16 fanout382 (.A(_05853_),
    .X(net382));
 sky130_fd_sc_hd__buf_12 fanout383 (.A(_05852_),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_16 fanout384 (.A(_05852_),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_16 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_16 fanout386 (.A(_05847_),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_16 fanout387 (.A(_05845_),
    .X(net387));
 sky130_fd_sc_hd__buf_12 fanout388 (.A(_05845_),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_16 fanout389 (.A(_05838_),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_16 fanout390 (.A(_05838_),
    .X(net390));
 sky130_fd_sc_hd__buf_12 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_12 fanout392 (.A(_02095_),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_16 fanout393 (.A(_02025_),
    .X(net393));
 sky130_fd_sc_hd__buf_12 fanout394 (.A(_02025_),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_16 fanout395 (.A(_02021_),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_16 fanout396 (.A(_02021_),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_16 fanout397 (.A(_02018_),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_16 fanout398 (.A(_02018_),
    .X(net398));
 sky130_fd_sc_hd__buf_12 fanout399 (.A(_02017_),
    .X(net399));
 sky130_fd_sc_hd__buf_4 fanout4 (.A(_06814_),
    .X(net3722));
 sky130_fd_sc_hd__clkbuf_16 fanout400 (.A(_02017_),
    .X(net400));
 sky130_fd_sc_hd__buf_12 fanout401 (.A(_02013_),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_16 fanout402 (.A(_02013_),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_8 fanout403 (.A(_01952_),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_8 fanout404 (.A(_01952_),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_16 fanout405 (.A(_01834_),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_16 fanout406 (.A(_01834_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_16 fanout407 (.A(_01833_),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_16 fanout408 (.A(_01833_),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_16 fanout409 (.A(_01831_),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_16 fanout410 (.A(_01831_),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_16 fanout411 (.A(_01828_),
    .X(net411));
 sky130_fd_sc_hd__buf_8 fanout412 (.A(_01828_),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_16 fanout413 (.A(_01822_),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_16 fanout414 (.A(_01822_),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_16 fanout415 (.A(_01743_),
    .X(net415));
 sky130_fd_sc_hd__buf_8 fanout416 (.A(_01743_),
    .X(net416));
 sky130_fd_sc_hd__buf_8 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_12 fanout418 (.A(_01742_),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_16 fanout419 (.A(_01741_),
    .X(net419));
 sky130_fd_sc_hd__buf_12 fanout420 (.A(_01741_),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_16 fanout421 (.A(_06809_),
    .X(net421));
 sky130_fd_sc_hd__buf_12 fanout422 (.A(_06809_),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_16 fanout423 (.A(_05854_),
    .X(net423));
 sky130_fd_sc_hd__buf_12 fanout424 (.A(_05854_),
    .X(net424));
 sky130_fd_sc_hd__buf_8 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_12 fanout426 (.A(_05851_),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_16 fanout427 (.A(_05850_),
    .X(net427));
 sky130_fd_sc_hd__buf_8 fanout428 (.A(_05850_),
    .X(net428));
 sky130_fd_sc_hd__buf_12 fanout429 (.A(_05849_),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_16 fanout430 (.A(_05849_),
    .X(net430));
 sky130_fd_sc_hd__buf_12 fanout431 (.A(_05848_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_16 fanout432 (.A(_05848_),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_16 fanout433 (.A(_02026_),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_16 fanout434 (.A(_02026_),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_16 fanout435 (.A(_02022_),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_16 fanout436 (.A(_02022_),
    .X(net436));
 sky130_fd_sc_hd__buf_12 fanout437 (.A(_02020_),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_16 fanout438 (.A(_02020_),
    .X(net438));
 sky130_fd_sc_hd__buf_12 fanout439 (.A(_02016_),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_16 fanout440 (.A(_02016_),
    .X(net440));
 sky130_fd_sc_hd__buf_4 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_4 fanout442 (.A(_02009_),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(_02009_),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(_02009_),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(net3415),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(_02009_),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(_02008_),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(_02008_),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(_02008_),
    .X(net451));
 sky130_fd_sc_hd__buf_4 fanout452 (.A(net454),
    .X(net452));
 sky130_fd_sc_hd__buf_2 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(_02008_),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_16 fanout455 (.A(_01824_),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_16 fanout456 (.A(_01824_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_4 fanout458 (.A(_05928_),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_4 fanout460 (.A(_05927_),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_8 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_8 fanout462 (.A(_05860_),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_16 fanout463 (.A(_01825_),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_16 fanout464 (.A(_01825_),
    .X(net464));
 sky130_fd_sc_hd__buf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_4 fanout466 (.A(_05894_),
    .X(net466));
 sky130_fd_sc_hd__buf_8 fanout467 (.A(_02101_),
    .X(net467));
 sky130_fd_sc_hd__buf_8 fanout468 (.A(_02100_),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(_02100_),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_4 fanout470 (.A(_05858_),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_4 fanout471 (.A(_05858_),
    .X(net471));
 sky130_fd_sc_hd__buf_4 fanout472 (.A(_02844_),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_4 fanout474 (.A(net476),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_8 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_4 fanout476 (.A(_01979_),
    .X(net476));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_8 fanout478 (.A(_01975_),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_8 fanout479 (.A(_01804_),
    .X(net479));
 sky130_fd_sc_hd__buf_6 fanout480 (.A(_01804_),
    .X(net480));
 sky130_fd_sc_hd__buf_8 fanout482 (.A(_02078_),
    .X(net482));
 sky130_fd_sc_hd__buf_8 fanout483 (.A(_02078_),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_16 fanout484 (.A(_02071_),
    .X(net484));
 sky130_fd_sc_hd__buf_8 fanout485 (.A(_02070_),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_4 fanout487 (.A(_05893_),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_4 fanout488 (.A(_05893_),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_4 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_4 fanout490 (.A(_01791_),
    .X(net490));
 sky130_fd_sc_hd__buf_8 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_8 fanout492 (.A(_01790_),
    .X(net492));
 sky130_fd_sc_hd__buf_8 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__buf_8 fanout494 (.A(_01790_),
    .X(net494));
 sky130_fd_sc_hd__buf_8 fanout495 (.A(net497),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_8 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_8 fanout497 (.A(_01789_),
    .X(net497));
 sky130_fd_sc_hd__buf_8 fanout498 (.A(_01789_),
    .X(net498));
 sky130_fd_sc_hd__buf_4 fanout499 (.A(_01789_),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout5 (.A(_06813_),
    .X(net3723));
 sky130_fd_sc_hd__buf_8 fanout500 (.A(_01789_),
    .X(net500));
 sky130_fd_sc_hd__buf_4 fanout501 (.A(_01789_),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_8 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__buf_6 fanout503 (.A(_01788_),
    .X(net503));
 sky130_fd_sc_hd__buf_6 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_6 fanout505 (.A(_01788_),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_16 fanout506 (.A(_01772_),
    .X(net506));
 sky130_fd_sc_hd__buf_8 fanout507 (.A(_01772_),
    .X(net507));
 sky130_fd_sc_hd__buf_6 fanout508 (.A(net510),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_8 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_4 fanout510 (.A(_01771_),
    .X(net510));
 sky130_fd_sc_hd__buf_6 fanout511 (.A(_01771_),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_4 fanout512 (.A(_01771_),
    .X(net512));
 sky130_fd_sc_hd__buf_6 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_6 fanout514 (.A(_01771_),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_8 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_6 fanout516 (.A(_01771_),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_8 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_8 fanout518 (.A(_00009_),
    .X(net518));
 sky130_fd_sc_hd__buf_6 fanout519 (.A(_00009_),
    .X(net519));
 sky130_fd_sc_hd__buf_6 fanout520 (.A(_00009_),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_8 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__buf_4 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__buf_6 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_8 fanout524 (.A(_00008_),
    .X(net524));
 sky130_fd_sc_hd__buf_6 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_8 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_4 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_8 fanout528 (.A(_00008_),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_8 fanout529 (.A(net533),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_8 fanout530 (.A(net533),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_8 fanout531 (.A(net533),
    .X(net531));
 sky130_fd_sc_hd__buf_4 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_8 fanout533 (.A(_00007_),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_8 fanout534 (.A(_00007_),
    .X(net534));
 sky130_fd_sc_hd__buf_6 fanout535 (.A(_00007_),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_8 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_6 fanout537 (.A(_00007_),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_8 fanout538 (.A(net542),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_8 fanout539 (.A(net542),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_8 fanout540 (.A(net542),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_8 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_8 fanout542 (.A(_00006_),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_8 fanout543 (.A(net546),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_8 fanout544 (.A(net546),
    .X(net544));
 sky130_fd_sc_hd__buf_4 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(_00006_),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_8 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_6 fanout548 (.A(net551),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_8 fanout549 (.A(net551),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_8 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_8 fanout551 (.A(_00006_),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_8 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_4 fanout553 (.A(_00006_),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_8 fanout554 (.A(net556),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_8 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_4 fanout556 (.A(_00006_),
    .X(net556));
 sky130_fd_sc_hd__buf_8 fanout557 (.A(net561),
    .X(net557));
 sky130_fd_sc_hd__buf_8 fanout558 (.A(net561),
    .X(net558));
 sky130_fd_sc_hd__buf_8 fanout559 (.A(net561),
    .X(net559));
 sky130_fd_sc_hd__buf_8 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_16 fanout561 (.A(net576),
    .X(net561));
 sky130_fd_sc_hd__buf_8 fanout562 (.A(net576),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_4 fanout563 (.A(net576),
    .X(net563));
 sky130_fd_sc_hd__buf_8 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__buf_8 fanout565 (.A(net576),
    .X(net565));
 sky130_fd_sc_hd__buf_8 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__buf_8 fanout567 (.A(net570),
    .X(net567));
 sky130_fd_sc_hd__buf_8 fanout568 (.A(net570),
    .X(net568));
 sky130_fd_sc_hd__buf_8 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_6 fanout570 (.A(net576),
    .X(net570));
 sky130_fd_sc_hd__buf_8 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_8 fanout572 (.A(net576),
    .X(net572));
 sky130_fd_sc_hd__buf_8 fanout573 (.A(net575),
    .X(net573));
 sky130_fd_sc_hd__buf_8 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_8 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__buf_8 fanout576 (.A(_00005_),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net3216),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_4 fanout578 (.A(net3216),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_8 fanout579 (.A(\dpath.alu.adder.in0[23] ),
    .X(net579));
 sky130_fd_sc_hd__buf_6 fanout580 (.A(\dpath.alu.adder.in0[22] ),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_8 fanout581 (.A(\dpath.alu.adder.in0[21] ),
    .X(net581));
 sky130_fd_sc_hd__buf_2 fanout582 (.A(\dpath.alu.adder.in0[21] ),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_8 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(\dpath.alu.adder.in0[20] ),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_8 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(\dpath.alu.adder.in0[19] ),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_8 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_8 fanout588 (.A(\dpath.alu.adder.in0[18] ),
    .X(net588));
 sky130_fd_sc_hd__buf_6 fanout589 (.A(net591),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_4 fanout591 (.A(\dpath.alu.adder.in0[17] ),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_8 fanout592 (.A(net594),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_8 fanout594 (.A(\dpath.alu.adder.in0[16] ),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_8 fanout595 (.A(net597),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_4 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_6 fanout597 (.A(\dpath.alu.adder.in0[15] ),
    .X(net597));
 sky130_fd_sc_hd__buf_4 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__buf_4 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_4 fanout6 (.A(_06813_),
    .X(net3724));
 sky130_fd_sc_hd__clkbuf_8 fanout600 (.A(\dpath.alu.adder.in0[14] ),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_8 fanout601 (.A(net603),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_4 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__buf_8 fanout603 (.A(\dpath.alu.adder.in0[13] ),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_8 fanout604 (.A(\dpath.alu.adder.in0[12] ),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_4 fanout605 (.A(\dpath.alu.adder.in0[12] ),
    .X(net605));
 sky130_fd_sc_hd__buf_6 fanout606 (.A(\dpath.alu.adder.in0[12] ),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_8 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__buf_8 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_8 fanout609 (.A(\dpath.alu.adder.in0[11] ),
    .X(net609));
 sky130_fd_sc_hd__buf_6 fanout610 (.A(\dpath.alu.adder.in0[10] ),
    .X(net610));
 sky130_fd_sc_hd__buf_6 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_8 fanout612 (.A(\dpath.alu.adder.in0[10] ),
    .X(net612));
 sky130_fd_sc_hd__buf_6 fanout613 (.A(net615),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_8 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_6 fanout615 (.A(\dpath.alu.adder.in0[9] ),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_8 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__buf_4 fanout617 (.A(\dpath.alu.adder.in0[8] ),
    .X(net617));
 sky130_fd_sc_hd__buf_6 fanout618 (.A(\dpath.alu.adder.in0[8] ),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 fanout619 (.A(\dpath.alu.adder.in0[8] ),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_8 fanout620 (.A(net623),
    .X(net620));
 sky130_fd_sc_hd__buf_4 fanout621 (.A(net623),
    .X(net621));
 sky130_fd_sc_hd__buf_6 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_8 fanout623 (.A(\dpath.alu.adder.in0[7] ),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_8 fanout624 (.A(net627),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout625 (.A(net627),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_8 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__buf_6 fanout627 (.A(\dpath.alu.adder.in0[6] ),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_8 fanout628 (.A(\dpath.alu.adder.in0[5] ),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_4 fanout629 (.A(\dpath.alu.adder.in0[5] ),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_8 fanout630 (.A(\dpath.alu.adder.in0[5] ),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_4 fanout631 (.A(\dpath.alu.adder.in0[5] ),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_8 fanout632 (.A(\dpath.alu.adder.in0[4] ),
    .X(net632));
 sky130_fd_sc_hd__buf_2 fanout633 (.A(\dpath.alu.adder.in0[4] ),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_8 fanout634 (.A(\dpath.alu.adder.in0[4] ),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_4 fanout635 (.A(\dpath.alu.adder.in0[4] ),
    .X(net635));
 sky130_fd_sc_hd__buf_4 fanout636 (.A(net638),
    .X(net636));
 sky130_fd_sc_hd__buf_2 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_4 fanout638 (.A(\dpath.alu.adder.in0[3] ),
    .X(net638));
 sky130_fd_sc_hd__buf_4 fanout639 (.A(net640),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_8 fanout640 (.A(\dpath.alu.adder.in0[3] ),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(net643),
    .X(net641));
 sky130_fd_sc_hd__buf_2 fanout642 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__buf_4 fanout643 (.A(\dpath.alu.adder.in0[2] ),
    .X(net643));
 sky130_fd_sc_hd__buf_4 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_8 fanout645 (.A(\dpath.alu.adder.in0[2] ),
    .X(net645));
 sky130_fd_sc_hd__buf_4 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_8 fanout647 (.A(\dpath.alu.adder.in0[1] ),
    .X(net647));
 sky130_fd_sc_hd__buf_4 fanout648 (.A(\dpath.alu.adder.in0[1] ),
    .X(net648));
 sky130_fd_sc_hd__buf_4 fanout649 (.A(\dpath.alu.adder.in0[1] ),
    .X(net649));
 sky130_fd_sc_hd__buf_4 fanout650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__buf_4 fanout651 (.A(\dpath.alu.adder.in0[0] ),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_8 fanout652 (.A(\dpath.alu.adder.in0[0] ),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_4 fanout653 (.A(\dpath.alu.adder.in0[0] ),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__buf_4 fanout655 (.A(\dpath.RF.wdata[31] ),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_4 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_4 fanout657 (.A(\dpath.RF.wdata[30] ),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_4 fanout658 (.A(net659),
    .X(net658));
 sky130_fd_sc_hd__buf_4 fanout659 (.A(net3689),
    .X(net659));
 sky130_fd_sc_hd__buf_4 fanout660 (.A(\dpath.RF.wdata[28] ),
    .X(net660));
 sky130_fd_sc_hd__buf_4 fanout661 (.A(net3637),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_4 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_4 fanout663 (.A(\dpath.RF.wdata[27] ),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_4 fanout664 (.A(\dpath.RF.wdata[26] ),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_4 fanout665 (.A(\dpath.RF.wdata[26] ),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 fanout666 (.A(net667),
    .X(net666));
 sky130_fd_sc_hd__buf_4 fanout667 (.A(\dpath.RF.wdata[25] ),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_4 fanout668 (.A(net670),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_2 fanout669 (.A(net670),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_4 fanout670 (.A(net3644),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_4 fanout671 (.A(net672),
    .X(net671));
 sky130_fd_sc_hd__buf_4 fanout672 (.A(\dpath.RF.wdata[23] ),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_4 fanout673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_4 fanout674 (.A(\dpath.RF.wdata[22] ),
    .X(net674));
 sky130_fd_sc_hd__buf_4 fanout675 (.A(net676),
    .X(net675));
 sky130_fd_sc_hd__buf_4 fanout676 (.A(net3623),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_4 fanout677 (.A(net679),
    .X(net677));
 sky130_fd_sc_hd__buf_2 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__buf_2 fanout679 (.A(net3630),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_4 fanout680 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_4 fanout681 (.A(net998),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_4 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_4 fanout683 (.A(\dpath.RF.wdata[18] ),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_4 fanout684 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__buf_4 fanout685 (.A(net1064),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__buf_4 fanout687 (.A(\dpath.RF.wdata[16] ),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_4 fanout689 (.A(\dpath.RF.wdata[15] ),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_4 fanout690 (.A(net691),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_4 fanout691 (.A(net3718),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_4 fanout692 (.A(\dpath.RF.wdata[13] ),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_4 fanout693 (.A(\dpath.RF.wdata[13] ),
    .X(net693));
 sky130_fd_sc_hd__buf_4 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__buf_4 fanout695 (.A(\dpath.RF.wdata[12] ),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_4 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__buf_4 fanout697 (.A(\dpath.RF.wdata[11] ),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_4 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__buf_4 fanout699 (.A(net1078),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_4 fanout700 (.A(net701),
    .X(net700));
 sky130_fd_sc_hd__buf_4 fanout701 (.A(\dpath.RF.wdata[9] ),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_4 fanout702 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__buf_4 fanout703 (.A(net1180),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_4 fanout704 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__buf_4 fanout705 (.A(\dpath.RF.wdata[7] ),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_4 fanout706 (.A(net707),
    .X(net706));
 sky130_fd_sc_hd__buf_4 fanout707 (.A(net1360),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_4 fanout708 (.A(net709),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_4 fanout709 (.A(\dpath.RF.wdata[5] ),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_4 fanout710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__buf_4 fanout711 (.A(\dpath.RF.wdata[4] ),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_4 fanout712 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__buf_4 fanout713 (.A(net3271),
    .X(net713));
 sky130_fd_sc_hd__buf_4 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__buf_4 fanout715 (.A(net1374),
    .X(net715));
 sky130_fd_sc_hd__buf_4 fanout716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__buf_4 fanout717 (.A(\dpath.RF.wdata[1] ),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_4 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__buf_4 fanout719 (.A(net3310),
    .X(net719));
 sky130_fd_sc_hd__buf_4 fanout720 (.A(\dpath.alu.adder.in1[24] ),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_8 fanout721 (.A(\dpath.alu.adder.in1[23] ),
    .X(net721));
 sky130_fd_sc_hd__buf_6 fanout722 (.A(\dpath.alu.adder.in1[22] ),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_8 fanout723 (.A(\dpath.alu.adder.in1[21] ),
    .X(net723));
 sky130_fd_sc_hd__buf_2 fanout724 (.A(\dpath.alu.adder.in1[21] ),
    .X(net724));
 sky130_fd_sc_hd__buf_6 fanout725 (.A(\dpath.alu.adder.in1[20] ),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_8 fanout726 (.A(\dpath.alu.adder.in1[19] ),
    .X(net726));
 sky130_fd_sc_hd__buf_4 fanout727 (.A(\dpath.alu.adder.in1[19] ),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_8 fanout728 (.A(net729),
    .X(net728));
 sky130_fd_sc_hd__buf_6 fanout729 (.A(\dpath.alu.adder.in1[18] ),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_8 fanout730 (.A(\dpath.alu.adder.in1[17] ),
    .X(net730));
 sky130_fd_sc_hd__buf_4 fanout731 (.A(\dpath.alu.adder.in1[17] ),
    .X(net731));
 sky130_fd_sc_hd__buf_4 fanout732 (.A(net733),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_8 fanout733 (.A(\dpath.alu.adder.in1[16] ),
    .X(net733));
 sky130_fd_sc_hd__buf_4 fanout734 (.A(net735),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_8 fanout735 (.A(\dpath.alu.adder.in1[15] ),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_8 fanout736 (.A(net738),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_4 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_8 fanout738 (.A(\dpath.alu.adder.in1[14] ),
    .X(net738));
 sky130_fd_sc_hd__buf_4 fanout739 (.A(\dpath.alu.adder.in1[13] ),
    .X(net739));
 sky130_fd_sc_hd__buf_4 fanout740 (.A(net742),
    .X(net740));
 sky130_fd_sc_hd__buf_2 fanout741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_4 fanout742 (.A(\dpath.alu.adder.in1[13] ),
    .X(net742));
 sky130_fd_sc_hd__buf_4 fanout743 (.A(\dpath.alu.adder.in1[12] ),
    .X(net743));
 sky130_fd_sc_hd__buf_4 fanout744 (.A(net746),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_4 fanout745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 fanout746 (.A(\dpath.alu.adder.in1[12] ),
    .X(net746));
 sky130_fd_sc_hd__buf_4 fanout747 (.A(\dpath.alu.adder.in1[11] ),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(net750),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_2 fanout750 (.A(\dpath.alu.adder.in1[11] ),
    .X(net750));
 sky130_fd_sc_hd__buf_4 fanout751 (.A(\dpath.alu.adder.in1[10] ),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(net753),
    .X(net752));
 sky130_fd_sc_hd__buf_4 fanout753 (.A(\dpath.alu.adder.in1[10] ),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(\dpath.alu.adder.in1[9] ),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_8 fanout755 (.A(\dpath.alu.adder.in1[9] ),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_8 fanout756 (.A(\dpath.alu.adder.in1[9] ),
    .X(net756));
 sky130_fd_sc_hd__buf_4 fanout757 (.A(\dpath.alu.adder.in1[8] ),
    .X(net757));
 sky130_fd_sc_hd__buf_4 fanout758 (.A(net759),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_8 fanout759 (.A(\dpath.alu.adder.in1[8] ),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_8 fanout760 (.A(net763),
    .X(net760));
 sky130_fd_sc_hd__buf_6 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_8 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_8 fanout763 (.A(\dpath.alu.adder.in1[7] ),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_8 fanout764 (.A(\dpath.alu.adder.in1[6] ),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_8 fanout765 (.A(net767),
    .X(net765));
 sky130_fd_sc_hd__buf_6 fanout766 (.A(net767),
    .X(net766));
 sky130_fd_sc_hd__buf_4 fanout767 (.A(\dpath.alu.adder.in1[6] ),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_8 fanout768 (.A(net771),
    .X(net768));
 sky130_fd_sc_hd__buf_6 fanout769 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_8 fanout770 (.A(net771),
    .X(net770));
 sky130_fd_sc_hd__buf_4 fanout771 (.A(\dpath.alu.adder.in1[5] ),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_8 fanout772 (.A(net775),
    .X(net772));
 sky130_fd_sc_hd__buf_4 fanout773 (.A(net775),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_8 fanout774 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_8 fanout775 (.A(\dpath.alu.adder.in1[4] ),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_8 fanout776 (.A(\dpath.alu.adder.in1[3] ),
    .X(net776));
 sky130_fd_sc_hd__buf_4 fanout777 (.A(\dpath.alu.adder.in1[3] ),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__buf_6 fanout779 (.A(\dpath.alu.adder.in1[3] ),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_8 fanout780 (.A(net782),
    .X(net780));
 sky130_fd_sc_hd__buf_4 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__buf_4 fanout782 (.A(\dpath.alu.adder.in1[2] ),
    .X(net782));
 sky130_fd_sc_hd__buf_4 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__buf_4 fanout784 (.A(\dpath.alu.adder.in1[1] ),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_8 fanout785 (.A(\dpath.alu.adder.in1[1] ),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_8 fanout786 (.A(\dpath.alu.adder.in1[0] ),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 fanout787 (.A(\dpath.alu.adder.in1[0] ),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_8 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_8 fanout789 (.A(\dpath.alu.adder.in1[0] ),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_8 fanout790 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__buf_6 fanout791 (.A(net3665),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_8 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_6 fanout793 (.A(net3677),
    .X(net793));
 sky130_fd_sc_hd__buf_8 fanout794 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__buf_8 fanout795 (.A(_00003_),
    .X(net795));
 sky130_fd_sc_hd__buf_6 fanout796 (.A(net797),
    .X(net796));
 sky130_fd_sc_hd__buf_8 fanout797 (.A(_00002_),
    .X(net797));
 sky130_fd_sc_hd__buf_6 fanout798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__buf_8 fanout799 (.A(_00002_),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_8 fanout800 (.A(net804),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_8 fanout801 (.A(net804),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_8 fanout802 (.A(net804),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_8 fanout803 (.A(net804),
    .X(net803));
 sky130_fd_sc_hd__buf_8 fanout804 (.A(net808),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_8 fanout805 (.A(net808),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_8 fanout806 (.A(net808),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_8 fanout807 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__buf_4 fanout808 (.A(_00001_),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_8 fanout809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_8 fanout810 (.A(_00001_),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_8 fanout811 (.A(net813),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_8 fanout812 (.A(net813),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_4 fanout813 (.A(_00001_),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_8 fanout814 (.A(_00001_),
    .X(net814));
 sky130_fd_sc_hd__buf_2 fanout815 (.A(_00001_),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_8 fanout816 (.A(net818),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_8 fanout817 (.A(net818),
    .X(net817));
 sky130_fd_sc_hd__buf_4 fanout818 (.A(_00001_),
    .X(net818));
 sky130_fd_sc_hd__buf_6 fanout819 (.A(net821),
    .X(net819));
 sky130_fd_sc_hd__buf_6 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__buf_6 fanout821 (.A(_00000_),
    .X(net821));
 sky130_fd_sc_hd__buf_8 fanout822 (.A(net824),
    .X(net822));
 sky130_fd_sc_hd__buf_8 fanout823 (.A(net824),
    .X(net823));
 sky130_fd_sc_hd__buf_6 fanout824 (.A(_00000_),
    .X(net824));
 sky130_fd_sc_hd__buf_6 fanout825 (.A(net829),
    .X(net825));
 sky130_fd_sc_hd__buf_6 fanout826 (.A(net828),
    .X(net826));
 sky130_fd_sc_hd__buf_6 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__buf_4 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_4 fanout829 (.A(_00000_),
    .X(net829));
 sky130_fd_sc_hd__buf_8 fanout830 (.A(net832),
    .X(net830));
 sky130_fd_sc_hd__buf_8 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_6 fanout832 (.A(net842),
    .X(net832));
 sky130_fd_sc_hd__buf_6 fanout833 (.A(net835),
    .X(net833));
 sky130_fd_sc_hd__buf_8 fanout834 (.A(net835),
    .X(net834));
 sky130_fd_sc_hd__buf_8 fanout835 (.A(net842),
    .X(net835));
 sky130_fd_sc_hd__buf_6 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__buf_6 fanout837 (.A(net842),
    .X(net837));
 sky130_fd_sc_hd__buf_6 fanout838 (.A(net842),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 fanout839 (.A(net842),
    .X(net839));
 sky130_fd_sc_hd__buf_6 fanout840 (.A(net842),
    .X(net840));
 sky130_fd_sc_hd__buf_4 fanout841 (.A(net842),
    .X(net841));
 sky130_fd_sc_hd__buf_6 fanout842 (.A(_00000_),
    .X(net842));
 sky130_fd_sc_hd__buf_4 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__buf_4 fanout844 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__buf_4 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout846 (.A(net850),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 fanout847 (.A(net849),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_4 fanout848 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_8 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_8 fanout850 (.A(net862),
    .X(net850));
 sky130_fd_sc_hd__buf_4 fanout851 (.A(net859),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_4 fanout852 (.A(net859),
    .X(net852));
 sky130_fd_sc_hd__buf_4 fanout853 (.A(net859),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 fanout854 (.A(net855),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_4 fanout855 (.A(net859),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 fanout856 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_2 fanout857 (.A(net859),
    .X(net857));
 sky130_fd_sc_hd__buf_4 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_4 fanout859 (.A(net861),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__buf_2 fanout861 (.A(net862),
    .X(net861));
 sky130_fd_sc_hd__buf_4 fanout862 (.A(_01792_),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_4 fanout863 (.A(net864),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_4 fanout864 (.A(net865),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_8 fanout865 (.A(net879),
    .X(net865));
 sky130_fd_sc_hd__buf_4 fanout866 (.A(net868),
    .X(net866));
 sky130_fd_sc_hd__buf_2 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_2 fanout868 (.A(net871),
    .X(net868));
 sky130_fd_sc_hd__buf_4 fanout869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_4 fanout870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__buf_2 fanout871 (.A(net872),
    .X(net871));
 sky130_fd_sc_hd__buf_4 fanout872 (.A(net879),
    .X(net872));
 sky130_fd_sc_hd__buf_4 fanout873 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__buf_2 fanout874 (.A(net876),
    .X(net874));
 sky130_fd_sc_hd__buf_4 fanout875 (.A(net876),
    .X(net875));
 sky130_fd_sc_hd__buf_4 fanout876 (.A(net879),
    .X(net876));
 sky130_fd_sc_hd__buf_2 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 fanout878 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__buf_6 fanout879 (.A(_01792_),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_8 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_8 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout882 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_8 fanout883 (.A(net889),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_8 fanout884 (.A(net889),
    .X(net884));
 sky130_fd_sc_hd__buf_4 fanout885 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_4 fanout886 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__buf_4 fanout887 (.A(net888),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_8 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_8 fanout889 (.A(net894),
    .X(net889));
 sky130_fd_sc_hd__buf_4 fanout890 (.A(net893),
    .X(net890));
 sky130_fd_sc_hd__buf_2 fanout891 (.A(net893),
    .X(net891));
 sky130_fd_sc_hd__buf_6 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_8 fanout893 (.A(net894),
    .X(net893));
 sky130_fd_sc_hd__buf_6 fanout894 (.A(net161),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\dpath.csrw_out_MW.d[13] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_01458_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_01467_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_00696_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\dpath.RF.R[7][29] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_00039_),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\dpath.RF.R[22][1] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_00351_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\dpath.RF.R[27][1] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_00962_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\dpath.RF.R[19][26] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_00344_),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\dpath.RF.R[9][12] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\dpath.csrw_out_MW.d[28] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_00717_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\dpath.RF.R[21][16] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_00430_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\dpath.RF.R[12][10] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_01580_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\dpath.RF.R[26][14] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_00911_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\dpath.RF.R[14][19] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_01300_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\dpath.RF.R[7][30] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_01213_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_00040_),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\dpath.RF.R[14][6] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_01287_),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\dpath.RF.R[12][6] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_01576_),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\dpath.RF.R[6][5] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_00047_),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\dpath.RF.R[19][3] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_00321_),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\dpath.RF.R[6][6] ),
    .X(net1924));
 sky130_fd_sc_hd__buf_1 hold103 (.A(\dpath.RF.wdata[19] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_00048_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\dpath.RF.R[14][10] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_01291_),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\dpath.RF.R[2][29] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_00830_),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\dpath.RF.R[7][16] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_00026_),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\dpath.RF.R[26][27] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_00924_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\dpath.RF.R[14][0] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_00433_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_01281_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\dpath.RF.R[26][19] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_00916_),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\dpath.RF.R[13][2] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_01475_),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\dpath.RF.R[4][22] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_00096_),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\dpath.RF.R[30][6] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_01645_),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\dpath.RF.R[21][10] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\ctrl.inst_X[24] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_00424_),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\dpath.RF.R[11][8] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_00937_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\dpath.RF.R[8][6] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_00999_),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\dpath.RF.R[5][18] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_00220_),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\dpath.RF.R[10][10] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_00843_),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\dpath.RF.R[28][17] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_00255_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_00882_),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\dpath.RF.R[17][17] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_00463_),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\dpath.RF.R[7][3] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_00013_),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\dpath.RF.R[22][13] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_00363_),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\dpath.RF.R[25][18] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_00755_),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\dpath.RF.R[23][13] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\dpath.csrw_out_DX.q[13] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_00681_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\dpath.RF.R[1][18] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_00528_),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\dpath.RF.R[3][14] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_00184_),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\dpath.csrw_out_DX.q[11] ),
    .X(net1970));
 sky130_fd_sc_hd__buf_1 hold1076 (.A(_01452_),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\dpath.RF.R[28][25] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_00890_),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\dpath.RF.R[18][28] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_01454_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_00634_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\dpath.RF.R[17][21] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_00467_),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\dpath.RF.R[19][16] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_00334_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\dpath.RF.R[8][20] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_01013_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\dpath.RF.R[11][29] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_00958_),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\dpath.RF.R[6][10] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\dpath.csrw_out_DX.q[27] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_00052_),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\dpath.RF.R[18][1] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_00607_),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\dpath.RF.R[19][7] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_00325_),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\dpath.RF.R[16][28] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_00570_),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\dpath.RF.R[14][4] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_01285_),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\dpath.RF.R[28][7] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\ctrl.inst_X[28] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_01468_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_00872_),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\dpath.RF.R[5][2] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_00204_),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\dpath.RF.R[8][3] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_00996_),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\dpath.RF.R[11][27] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_00956_),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\dpath.RF.R[4][8] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_00082_),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\dpath.RF.R[16][12] ),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\ctrl.inst_M[24] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_00554_),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\dpath.RF.R[8][18] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_01011_),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\dpath.RF.R[19][5] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_00323_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\dpath.RF.R[22][16] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_00366_),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\dpath.RF.R[11][13] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_00942_),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\dpath.RF.R[30][21] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_00310_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_01660_),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\dpath.RF.R[15][9] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_00583_),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\dpath.RF.R[2][23] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_00824_),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\dpath.RF.R[1][16] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_00526_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\dpath.RF.R[18][21] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_00627_),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\dpath.RF.R[15][30] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\dpath.csrw_out_DX.q[30] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_00604_),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\dpath.RF.R[1][8] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_00518_),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\dpath.RF.R[30][13] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_01652_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\dpath.RF.R[5][24] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_00226_),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\dpath.RF.R[27][8] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_00969_),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\dpath.RF.R[6][28] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_01471_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_00070_),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\dpath.RF.R[23][5] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_00673_),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\dpath.RF.R[21][13] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_00427_),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\dpath.RF.R[13][29] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_01502_),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\dpath.RF.R[5][31] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_00233_),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\dpath.RF.R[25][24] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\dpath.csrw_out_MW.d[4] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_00761_),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\dpath.RF.R[10][13] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_00846_),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\dpath.RF.R[5][4] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_00206_),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\dpath.RF.R[12][3] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_01573_),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\dpath.RF.R[23][15] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_00683_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\dpath.RF.R[27][16] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_01189_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_00977_),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\dpath.RF.R[20][9] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_00487_),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\dpath.RF.R[24][2] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_01604_),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\ctrl.d2c_inst[0] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_00264_),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\dpath.RF.R[27][5] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_00966_),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\dpath.RF.R[19][18] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\dpath.csrw_out_MW.d[23] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_00336_),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\dpath.RF.R[14][21] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_01302_),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\dpath.RF.R[27][20] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_00981_),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\dpath.RF.R[12][2] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_01572_),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\dpath.RF.R[3][27] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_00197_),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\dpath.RF.R[27][2] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_01208_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_00963_),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\dpath.RF.R[20][4] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_00482_),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\dpath.RF.R[21][0] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_00414_),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\dpath.RF.R[8][26] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_01019_),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\dpath.RF.R[23][29] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_00697_),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\dpath.RF.R[2][11] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\dpath.sd_DX.q[17] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_00812_),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\dpath.RF.R[2][10] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_00811_),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\dpath.RF.R[28][20] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_00885_),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\dpath.RF.R[2][12] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_00813_),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\dpath.csrw_out_DX.q[5] ),
    .X(net2092));
 sky130_fd_sc_hd__buf_1 hold1198 (.A(_01446_),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\dpath.RF.R[4][13] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00259_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_00399_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_00087_),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\dpath.RF.R[23][0] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_00668_),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\dpath.RF.R[21][17] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_00431_),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\dpath.RF.R[9][14] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_00719_),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\dpath.RF.R[7][9] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_00019_),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\dpath.RF.R[15][3] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\dpath.csrw_out_DX.q[16] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_00577_),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\dpath.RF.R[20][19] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_00497_),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\dpath.RF.R[15][19] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_00593_),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\dpath.RF.R[26][5] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_00902_),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\dpath.RF.R[27][29] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_00990_),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\dpath.RF.R[1][31] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_01457_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_00541_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\dpath.RF.R[24][17] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_01619_),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\dpath.RF.R[23][10] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_00678_),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\dpath.RF.R[9][22] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_00727_),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\dpath.RF.R[10][12] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_00845_),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\dpath.RF.R[1][30] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\dpath.csrw_out_DX.q[10] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_00540_),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\dpath.RF.R[8][23] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_01016_),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\dpath.RF.R[22][7] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_00357_),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\dpath.RF.R[22][31] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_00381_),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\dpath.RF.R[7][19] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_00029_),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\dpath.RF.R[19][29] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_01451_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_00347_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\dpath.RF.R[11][24] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_00953_),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\dpath.RF.R[26][21] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_00918_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\dpath.RF.R[2][26] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_00827_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\dpath.RF.R[28][15] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_00880_),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\dpath.RF.R[28][11] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\dpath.sd_DX.q[15] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_00876_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\dpath.RF.R[20][23] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_00501_),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\dpath.RF.R[26][2] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_00899_),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\dpath.RF.R[24][31] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_01633_),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\dpath.RF.R[10][18] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_00851_),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\dpath.RF.R[14][15] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_00397_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_01296_),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\dpath.RF.R[7][17] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_00027_),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\dpath.RF.R[16][0] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_00542_),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\dpath.RF.R[20][17] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_00495_),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\dpath.RF.R[26][24] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_00921_),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\dpath.RF.R[30][9] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\ctrl.inst_M[0] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_01648_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\dpath.RF.R[23][31] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_00699_),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\dpath.RF.R[20][13] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_00491_),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\dpath.RF.R[24][1] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(_01603_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\dpath.RF.R[6][22] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(_00064_),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\dpath.RF.R[15][31] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_00291_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(_00605_),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\dpath.RF.R[1][4] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_00514_),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\dpath.RF.R[13][14] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_01487_),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\dpath.RF.R[1][14] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_00524_),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\dpath.RF.R[4][19] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_00093_),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\dpath.RF.R[26][6] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\dpath.sd_DX.q[12] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_00903_),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\dpath.RF.R[18][5] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(_00611_),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\dpath.RF.R[21][23] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(_00437_),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\dpath.RF.R[17][24] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(_00470_),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\dpath.RF.R[27][14] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_00975_),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\dpath.RF.R[29][22] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\dpath.sd_DX.q[1] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_00394_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(_00160_),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\dpath.RF.R[6][16] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_00058_),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\dpath.RF.R[28][9] ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_00874_),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\dpath.RF.R[7][12] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(_00022_),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\dpath.RF.R[8][17] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(_01010_),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\dpath.RF.R[27][3] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\dpath.sd_DX.q[9] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(_00964_),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\dpath.RF.R[20][25] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_00503_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\dpath.RF.R[13][16] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(_01489_),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\dpath.RF.R[7][13] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_00023_),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\dpath.RF.R[2][8] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(_00809_),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\dpath.RF.R[3][15] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_00391_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(_00185_),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\dpath.RF.R[13][21] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(_01494_),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\dpath.RF.R[24][8] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_01610_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\dpath.RF.R[18][2] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(_00608_),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\dpath.RF.R[12][25] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_01595_),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\dpath.RF.R[7][14] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\dpath.csrw_out_DX.q[23] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(_00024_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\dpath.RF.R[12][29] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(_01599_),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\dpath.RF.R[24][3] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_01605_),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\dpath.RF.R[28][18] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_00883_),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\dpath.RF.R[4][27] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(_00101_),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\dpath.RF.R[6][24] ),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_01464_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(_00066_),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\dpath.RF.R[2][5] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(_00806_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\dpath.RF.R[29][31] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(_00169_),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\dpath.RF.R[15][29] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_00603_),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\dpath.RF.R[16][14] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_00556_),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\dpath.RF.R[4][28] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\dpath.sd_DX.q[11] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(_00102_),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\dpath.RF.R[8][5] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(_00998_),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\dpath.RF.R[11][5] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(_00934_),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\dpath.RF.R[13][1] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(_01474_),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\dpath.RF.R[7][6] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_00016_),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\dpath.RF.R[15][2] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_00393_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_00576_),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\dpath.RF.R[3][12] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_00182_),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\dpath.RF.R[27][22] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_00983_),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\dpath.RF.R[12][27] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_01597_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\dpath.RF.R[17][7] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_00453_),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\dpath.RF.R[16][23] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\dpath.csrw_out_MW.d[20] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(_00565_),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\dpath.RF.R[15][14] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_00588_),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\dpath.RF.R[15][17] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_00591_),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\dpath.RF.R[9][10] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(_00715_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\dpath.RF.R[8][12] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_01005_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\dpath.RF.R[26][0] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_01205_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(_00897_),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\dpath.RF.R[4][21] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(_00095_),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\dpath.RF.R[10][16] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_00849_),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\dpath.RF.R[26][11] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_00908_),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\dpath.RF.R[4][20] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(_00094_),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\dpath.RF.R[27][31] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\dpath.sd_DX.q[19] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_00992_),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\dpath.RF.R[17][9] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(_00455_),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\dpath.RF.R[23][30] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(_00698_),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\dpath.RF.R[30][14] ),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(_01653_),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\dpath.RF.R[2][17] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_00818_),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\dpath.RF.R[11][4] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00383_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_00401_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(_00933_),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\dpath.RF.R[2][2] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(_00803_),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\dpath.RF.R[3][28] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_00198_),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\dpath.RF.R[13][19] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_01492_),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\dpath.RF.R[11][15] ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_00944_),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\dpath.RF.R[7][31] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\dpath.csrw_out_MW.d[29] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_00041_),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\dpath.RF.R[25][21] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_00758_),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\dpath.RF.R[9][16] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_00721_),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\dpath.RF.R[18][16] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_00622_),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\dpath.RF.R[13][8] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(_01481_),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\dpath.RF.R[17][23] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_01214_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(_00469_),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\dpath.RF.R[4][10] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_00084_),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\dpath.RF.R[21][20] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(_00434_),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\dpath.RF.R[6][3] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(_00045_),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\dpath.RF.R[19][4] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(_00322_),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\dpath.RF.R[20][30] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\dpath.sd_DX.q[14] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_00508_),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\dpath.RF.R[28][16] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(_00881_),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\dpath.RF.R[17][19] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(_00465_),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\dpath.RF.R[5][19] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_00221_),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\dpath.RF.R[2][15] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(_00816_),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\dpath.RF.R[27][21] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_00396_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_00982_),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\dpath.RF.R[17][30] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(_00476_),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\dpath.RF.R[5][16] ),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(_00218_),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\dpath.RF.R[27][6] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(_00967_),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\dpath.RF.R[9][18] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_00723_),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\dpath.RF.R[1][15] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\ctrl.inst_M[25] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(_00525_),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\dpath.RF.R[5][29] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(_00231_),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\dpath.RF.R[19][9] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_00327_),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\dpath.RF.R[16][25] ),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_00567_),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\dpath.RF.R[21][25] ),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(_00439_),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\dpath.RF.R[3][7] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_00311_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(_00177_),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\dpath.RF.R[25][20] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(_00757_),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\dpath.RF.R[16][31] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(_00573_),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\dpath.RF.R[21][31] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(_00445_),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\dpath.RF.R[21][15] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(_00429_),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\dpath.RF.R[24][24] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\dpath.csrw_out_MW.d[12] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(_01626_),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\dpath.RF.R[8][8] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_01001_),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\dpath.RF.R[14][5] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_01286_),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\dpath.RF.R[19][25] ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(_00343_),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\dpath.RF.R[11][7] ),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(_00936_),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\dpath.RF.R[29][30] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_01197_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(_00168_),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\dpath.RF.R[7][24] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(_00034_),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\dpath.RF.R[9][21] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(_00726_),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\dpath.RF.R[21][4] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(_00418_),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\dpath.RF.R[25][23] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(_00760_),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\dpath.RF.R[4][5] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\dpath.sd_DX.q[13] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_00079_),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\dpath.RF.R[25][28] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(_00765_),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\dpath.RF.R[10][5] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(_00838_),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\dpath.RF.R[7][21] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(_00031_),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\dpath.RF.R[30][1] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(_01640_),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\dpath.RF.R[1][13] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\ctrl.inst_X[27] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_00395_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(_00523_),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\dpath.RF.R[25][13] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(_00750_),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\dpath.RF.R[5][25] ),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(_00227_),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\dpath.RF.R[2][21] ),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(_00822_),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\dpath.RF.R[3][30] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_00200_),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\dpath.RF.R[13][17] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\dpath.sd_DX.q[8] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(_01490_),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\ctrl.d2c_inst[1] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(_00265_),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\dpath.RF.R[23][27] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(_00695_),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\dpath.RF.R[10][7] ),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(_00840_),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\dpath.RF.R[17][4] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(_00450_),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\dpath.RF.R[12][12] ),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_00390_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(_01582_),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(\dpath.RF.R[27][9] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(_00970_),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\dpath.RF.R[3][10] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(_00180_),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\dpath.RF.R[3][3] ),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(_00173_),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\dpath.RF.R[19][12] ),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(_00330_),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\dpath.RF.R[24][5] ),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\dpath.csrw_out_MW.d[24] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(_01607_),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\dpath.RF.R[19][6] ),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_00324_),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\dpath.RF.R[26][26] ),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_00923_),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\dpath.RF.R[15][28] ),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(_00602_),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\dpath.RF.R[7][10] ),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_00020_),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\dpath.RF.R[26][17] ),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_01209_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(_00914_),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\dpath.RF.R[14][14] ),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(_01295_),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\dpath.RF.R[30][8] ),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_01647_),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\dpath.RF.R[2][7] ),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(_00808_),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\dpath.RF.R[3][2] ),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_00172_),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\dpath.RF.R[31][16] ),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\dpath.sd_DX.q[23] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(_00122_),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\dpath.RF.R[7][15] ),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(_00025_),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\dpath.RF.R[16][19] ),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_00561_),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\dpath.RF.R[23][14] ),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(_00682_),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\dpath.RF.R[10][19] ),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(_00852_),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\dpath.RF.R[20][6] ),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_00405_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_00484_),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\dpath.RF.R[16][24] ),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(_00566_),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\dpath.RF.R[31][4] ),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(_00110_),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\dpath.RF.R[23][19] ),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_00687_),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\dpath.RF.R[23][8] ),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_00676_),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\dpath.RF.R[6][14] ),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\dpath.RF.R[0][27] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(_00056_),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\dpath.RF.R[29][26] ),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_00164_),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\dpath.RF.R[25][15] ),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(_00752_),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\dpath.RF.R[8][4] ),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_00997_),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\dpath.RF.R[8][21] ),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_01014_),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\dpath.RF.R[2][9] ),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_00796_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(_00810_),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\dpath.RF.R[8][16] ),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_01009_),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\dpath.RF.R[8][10] ),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(_01003_),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\dpath.RF.R[11][9] ),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(_00938_),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\dpath.RF.R[1][5] ),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_00515_),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\dpath.RF.R[2][14] ),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\dpath.csrw_out_MW.d[1] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(_00815_),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\dpath.RF.R[31][1] ),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(_00107_),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\dpath.RF.R[15][13] ),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(_00587_),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\dpath.RF.R[23][25] ),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(_00693_),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\dpath.RF.R[21][27] ),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(_00441_),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\dpath.RF.R[22][26] ),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00258_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_01186_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_00376_),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\dpath.RF.R[12][28] ),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_01598_),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\dpath.RF.R[11][0] ),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_00929_),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\dpath.RF.R[8][11] ),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_01004_),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\dpath.RF.R[24][18] ),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(_01620_),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\dpath.RF.R[13][27] ),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\dpath.sd_DX.q[24] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(_01500_),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\dpath.RF.R[13][20] ),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_01493_),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\dpath.RF.R[3][13] ),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_00183_),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\dpath.RF.R[3][31] ),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(_00201_),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\dpath.RF.R[28][4] ),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(_00869_),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\dpath.RF.R[16][18] ),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_00406_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_00560_),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\dpath.RF.R[21][26] ),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(_00440_),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\dpath.RF.R[23][16] ),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_00684_),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\dpath.RF.R[19][28] ),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(_00346_),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\dpath.RF.R[3][17] ),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(_00187_),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\dpath.RF.R[27][28] ),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\dpath.RF.R[0][25] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(_00989_),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\dpath.RF.R[23][4] ),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_00672_),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\dpath.RF.R[25][19] ),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(_00756_),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\dpath.RF.R[11][14] ),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(_00943_),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\dpath.RF.R[21][2] ),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_00416_),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\dpath.RF.R[3][24] ),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_00794_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_00194_),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\dpath.RF.R[25][31] ),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(_00768_),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\dpath.RF.R[24][4] ),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_01606_),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\dpath.RF.R[22][11] ),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(_00361_),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\dpath.RF.R[5][1] ),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_00203_),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\dpath.RF.R[1][21] ),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\dpath.RF.R[0][0] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(_00531_),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\dpath.RF.R[9][11] ),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(_00716_),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\dpath.RF.R[4][1] ),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(_00075_),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\dpath.RF.R[30][7] ),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(_01646_),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\dpath.RF.R[6][26] ),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(_00068_),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\dpath.RF.R[24][27] ),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_00769_),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(_01629_),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\dpath.RF.R[30][0] ),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(_01639_),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\dpath.RF.R[3][22] ),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(_00192_),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\dpath.RF.R[21][11] ),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_00425_),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\dpath.RF.R[31][18] ),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_00124_),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\dpath.RF.R[30][3] ),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\dpath.sd_DX.q[25] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_01642_),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\dpath.RF.R[19][22] ),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(_00340_),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\dpath.RF.R[28][26] ),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_00891_),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\dpath.RF.R[16][17] ),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(_00559_),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\dpath.RF.R[29][24] ),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(_00162_),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\dpath.RF.R[22][5] ),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_00407_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_00355_),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\dpath.RF.R[31][15] ),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(_00121_),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\dpath.RF.R[19][24] ),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(_00342_),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\dpath.RF.R[10][15] ),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(_00848_),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\dpath.RF.R[6][27] ),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(_00069_),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\dpath.RF.R[7][5] ),
    .X(net2584));
 sky130_fd_sc_hd__buf_1 hold169 (.A(\dpath.RF.wdata[17] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(_00015_),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\dpath.RF.R[1][9] ),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(_00519_),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\dpath.RF.R[19][17] ),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(_00335_),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\dpath.RF.R[21][5] ),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(_00419_),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\dpath.RF.R[10][11] ),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_00844_),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\dpath.RF.R[31][21] ),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\ctrl.inst_X[30] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_00367_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(_00127_),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\dpath.RF.R[6][9] ),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(_00051_),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\dpath.RF.R[21][21] ),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(_00435_),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\dpath.RF.R[5][9] ),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(_00211_),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\dpath.RF.R[17][18] ),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(_00464_),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\dpath.RF.R[15][11] ),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\dpath.csrw_out_MW.d[30] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(_00585_),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\dpath.RF.R[29][6] ),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(_00144_),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\dpath.RF.R[15][6] ),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(_00580_),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\dpath.RF.R[27][23] ),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(_00984_),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\dpath.RF.R[29][1] ),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_00139_),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\dpath.RF.R[24][20] ),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_01215_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(_01622_),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\dpath.RF.R[29][25] ),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(_00163_),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\dpath.RF.R[4][17] ),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(_00091_),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\dpath.csrw_out_DX.q[1] ),
    .X(net2620));
 sky130_fd_sc_hd__buf_1 hold1726 (.A(_01442_),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\dpath.RF.R[19][13] ),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(_00331_),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\dpath.RF.R[31][10] ),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\dpath.sd_DX.q[0] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(_00116_),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\dpath.RF.R[13][23] ),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(_01496_),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\dpath.RF.R[29][4] ),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(_00142_),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(\dpath.RF.R[18][6] ),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(_00612_),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\dpath.RF.R[11][20] ),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(_00949_),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\dpath.RF.R[21][3] ),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_00382_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(_00417_),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\dpath.RF.R[29][29] ),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(_00167_),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\dpath.RF.R[31][23] ),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(_00129_),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\dpath.RF.R[4][15] ),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(_00089_),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\dpath.RF.R[19][19] ),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(_00337_),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\dpath.RF.R[3][8] ),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\dpath.sd_DX.q[6] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(_00178_),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\dpath.RF.R[4][4] ),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(_00078_),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\dpath.RF.R[9][2] ),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(_00707_),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\dpath.RF.R[26][13] ),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(_00910_),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\dpath.RF.R[14][23] ),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(_01304_),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\dpath.RF.R[7][0] ),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_00388_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(_00010_),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\dpath.RF.R[7][22] ),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(_00032_),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\dpath.RF.R[23][20] ),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(_00688_),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\dpath.RF.R[24][29] ),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(_01631_),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\dpath.RF.R[24][0] ),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(_01602_),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\dpath.RF.R[6][15] ),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\dpath.sd_DX.q[16] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(_00057_),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\dpath.RF.R[9][17] ),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(_00722_),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\dpath.RF.R[28][27] ),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(_00892_),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\dpath.RF.R[3][21] ),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(_00191_),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\dpath.RF.R[23][21] ),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(_00689_),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\dpath.RF.R[3][26] ),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_00398_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(_00196_),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\dpath.RF.R[15][26] ),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(_00600_),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\dpath.RF.R[15][15] ),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(_00589_),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\dpath.RF.R[25][8] ),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(_00745_),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\dpath.RF.R[28][8] ),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(_00873_),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\dpath.RF.R[4][16] ),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\dpath.RF.R[0][7] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_00090_),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\dpath.RF.R[17][31] ),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(_00477_),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\dpath.RF.R[31][17] ),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(_00123_),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\dpath.RF.R[27][7] ),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(_00968_),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\dpath.RF.R[8][1] ),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(_00994_),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\dpath.RF.R[27][15] ),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_00261_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_00776_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(_00976_),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\dpath.RF.R[7][18] ),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(_00028_),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\dpath.RF.R[23][12] ),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(_00680_),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\dpath.RF.R[29][5] ),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(_00143_),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\dpath.RF.R[31][29] ),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(_00135_),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\dpath.RF.R[10][26] ),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\dpath.sd_DX.q[20] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(_00859_),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\dpath.RF.R[19][14] ),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(_00332_),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\dpath.RF.R[24][21] ),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(_01623_),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\dpath.RF.R[29][20] ),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(_00158_),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\dpath.RF.R[4][31] ),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(_00105_),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\dpath.RF.R[17][12] ),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_00402_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(_00458_),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\dpath.RF.R[20][16] ),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(_00494_),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\dpath.RF.R[4][11] ),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(_00085_),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\dpath.RF.R[5][10] ),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(_00212_),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(\dpath.RF.R[22][8] ),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(_00358_),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(\dpath.RF.R[15][12] ),
    .X(net2724));
 sky130_fd_sc_hd__buf_1 hold183 (.A(\dpath.RF.wdata[10] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(_00586_),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(\dpath.RF.R[17][3] ),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(_00449_),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(\dpath.RF.R[18][14] ),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(_00620_),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\dpath.RF.R[17][13] ),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(_00459_),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\dpath.RF.R[20][26] ),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(_00504_),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\dpath.RF.R[4][9] ),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_00971_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(_00083_),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\dpath.RF.R[9][6] ),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(_00711_),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\dpath.RF.R[24][13] ),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(_01615_),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\dpath.RF.R[13][12] ),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(_01485_),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(\dpath.RF.R[3][18] ),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(_00188_),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\dpath.RF.R[31][0] ),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\dpath.RF.R[0][4] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(_00106_),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(\dpath.RF.R[19][11] ),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(_00329_),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(\dpath.RF.R[5][14] ),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(_00216_),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(\dpath.RF.R[3][23] ),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(_00193_),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(\dpath.RF.R[8][24] ),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(_01017_),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(\dpath.RF.R[4][14] ),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_00773_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(_00088_),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(\dpath.RF.R[20][27] ),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(_00505_),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(\dpath.RF.R[19][21] ),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(_00339_),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(\dpath.RF.R[18][12] ),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(_00618_),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(\dpath.RF.R[12][18] ),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(_01588_),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(\dpath.RF.R[4][30] ),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\dpath.RF.R[0][6] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(_00104_),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(\dpath.RF.R[1][20] ),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(_00530_),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(\dpath.RF.R[3][25] ),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(_00195_),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(\dpath.RF.R[31][20] ),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(_00126_),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(\dpath.RF.R[25][22] ),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(_00759_),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(\dpath.RF.R[6][12] ),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_00775_),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(_00054_),
    .X(net2775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\dpath.RF.R[27][4] ),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(_00965_),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(\dpath.RF.R[1][27] ),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(_00537_),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(\dpath.RF.R[13][6] ),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(_01479_),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\dpath.RF.R[5][6] ),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(_00208_),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(\dpath.RF.R[4][7] ),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\dpath.sd_DX.q[2] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(_00081_),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(\dpath.RF.R[2][0] ),
    .X(net2786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(_00801_),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(\dpath.RF.R[4][24] ),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(_00098_),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(\dpath.RF.R[25][30] ),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(_00767_),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(\dpath.RF.R[11][25] ),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(_00954_),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(\dpath.RF.R[3][11] ),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ctrl.inst_X[29] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_00384_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(_00181_),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(\dpath.RF.R[3][9] ),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(_00179_),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\dpath.RF.R[11][26] ),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(_00955_),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(\dpath.RF.R[21][18] ),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(_00432_),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(\dpath.RF.R[19][30] ),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(_00348_),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(\dpath.RF.R[2][20] ),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\dpath.sd_DX.q[18] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(_00821_),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(\dpath.RF.R[9][24] ),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(_00729_),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(\dpath.RF.R[4][29] ),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(_00103_),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(\dpath.RF.R[26][12] ),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(_00909_),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(\dpath.RF.R[11][17] ),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(_00946_),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(\dpath.RF.R[3][4] ),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_00400_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(_00174_),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(\dpath.RF.R[19][31] ),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(_00349_),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(\dpath.RF.R[25][16] ),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(_00753_),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(\dpath.RF.R[17][14] ),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(_00460_),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(\dpath.RF.R[23][24] ),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(_00692_),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(\dpath.RF.R[22][9] ),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\dpath.sd_DX.q[22] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(_00359_),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\dpath.RF.R[3][29] ),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(_00199_),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(\dpath.RF.R[21][12] ),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(_00426_),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(\dpath.RF.R[7][8] ),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(_00018_),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(\dpath.RF.R[13][7] ),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(_01480_),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(\dpath.RF.R[8][7] ),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_00404_),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(_01000_),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(\dpath.RF.R[31][19] ),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(_00125_),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(\dpath.RF.R[3][1] ),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(_00171_),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\dpath.RF.R[8][2] ),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(_00995_),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(\dpath.RF.R[30][22] ),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(_01661_),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(\dpath.RF.R[2][6] ),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\ctrl.inst_X[31] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(_00807_),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\dpath.RF.R[11][19] ),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(_00948_),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(\dpath.RF.R[7][28] ),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(_00038_),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(\dpath.RF.R[10][1] ),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(_00834_),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(\dpath.RF.R[29][28] ),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(_00166_),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(\dpath.RF.R[23][7] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_00262_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(_00675_),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(\dpath.RF.R[27][12] ),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(_00973_),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(\dpath.RF.R[15][21] ),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(_00595_),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(\dpath.RF.R[29][23] ),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(_00161_),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(\dpath.RF.R[15][27] ),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(_00601_),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(\dpath.RF.R[6][0] ),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\ctrl.inst_X[25] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(_00042_),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(\dpath.RF.R[5][13] ),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(_00215_),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(\ctrl.inst_X[13] ),
    .X(net2868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(_00249_),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(\dpath.RF.R[15][24] ),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(_00598_),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(\dpath.RF.R[15][25] ),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(_00599_),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(\dpath.RF.R[29][9] ),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_00256_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(_00147_),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(\dpath.RF.R[23][3] ),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(_00671_),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(\dpath.RF.R[25][10] ),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(_00747_),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(\dpath.RF.R[15][7] ),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(_00581_),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(\dpath.RF.R[15][23] ),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(_00597_),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(\dpath.RF.R[25][1] ),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\dpath.RF.R[24][10] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(_00738_),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(\dpath.RF.R[17][5] ),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(_00451_),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\dpath.RF.R[11][6] ),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(_00935_),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(\dpath.RF.R[20][31] ),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(_00509_),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(\dpath.RF.R[4][6] ),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(_00080_),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(\dpath.RF.R[6][17] ),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_01198_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00260_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_01612_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(_00059_),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(\dpath.RF.R[3][19] ),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(_00189_),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(\dpath.RF.R[31][31] ),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(_00137_),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(\dpath.RF.R[29][3] ),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(_00141_),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(\dpath.RF.R[25][6] ),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(_00743_),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(\dpath.RF.R[11][28] ),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\dpath.RF.R[0][21] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(_00957_),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(\dpath.RF.R[13][4] ),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(_01477_),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(\dpath.RF.R[15][5] ),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(_00579_),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(\dpath.RF.R[12][23] ),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(_01593_),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(\dpath.RF.R[11][2] ),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(_00931_),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(\dpath.RF.R[29][15] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00790_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(_00153_),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(\dpath.RF.R[6][13] ),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(_00055_),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(\dpath.RF.R[9][7] ),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(_00712_),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(\dpath.RF.R[29][8] ),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(_00146_),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(\dpath.RF.R[13][9] ),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(_01482_),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(\dpath.RF.R[17][0] ),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\dpath.RF.R[0][3] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(_00446_),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(\dpath.RF.R[7][20] ),
    .X(net2926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(_00030_),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(\dpath.RF.R[30][11] ),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(_01650_),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(\dpath.RF.R[27][26] ),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(_00987_),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(\dpath.RF.R[5][0] ),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(_00202_),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(\dpath.RF.R[20][7] ),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_00772_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(_00485_),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(\dpath.RF.R[15][22] ),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(_00596_),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(\dpath.RF.R[19][23] ),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(_00341_),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(\dpath.RF.R[6][30] ),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(_00072_),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(\dpath.RF.R[11][18] ),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(_00947_),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(\dpath.RF.R[4][2] ),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\dpath.RF.R[0][22] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(_00076_),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(\dpath.RF.R[15][16] ),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2052 (.A(_00590_),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(\dpath.RF.R[14][7] ),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(_01288_),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(\ctrl.inst_M[11] ),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(_01784_),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(\dpath.RF.R[31][7] ),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(_00113_),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(\dpath.RF.R[31][13] ),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_00791_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2060 (.A(_00119_),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(\dpath.RF.R[11][22] ),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2062 (.A(_00951_),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(\dpath.RF.R[31][9] ),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(_00115_),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(\dpath.RF.R[10][22] ),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2066 (.A(_00855_),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(\dpath.RF.R[9][1] ),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(_00706_),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(\dpath.RF.R[21][14] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\dpath.RF.R[0][20] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(_00428_),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2071 (.A(\dpath.RF.R[7][11] ),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(_00021_),
    .X(net2967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(\dpath.RF.R[13][25] ),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(_01498_),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(\dpath.RF.R[29][10] ),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2076 (.A(_00148_),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2077 (.A(\ctrl.inst_X[14] ),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(_00250_),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(\dpath.RF.R[3][16] ),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_00789_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(_00186_),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2081 (.A(\dpath.RF.R[31][14] ),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(_00120_),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(\dpath.RF.R[29][19] ),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(_00157_),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(\dpath.RF.R[17][1] ),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(_00447_),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2087 (.A(\dpath.RF.R[11][12] ),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2088 (.A(_00941_),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(\dpath.RF.R[29][21] ),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\dpath.sd_DX.q[21] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(_00159_),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(\dpath.RF.R[4][18] ),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(_00092_),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(\dpath.RF.R[21][6] ),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(_00420_),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(\dpath.RF.R[31][12] ),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(_00118_),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2097 (.A(\dpath.RF.R[14][12] ),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(_01293_),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(\dpath.RF.R[9][9] ),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\dpath.csrw_out_MW.d[8] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_00403_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(_00714_),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2101 (.A(\dpath.RF.R[27][17] ),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(_00978_),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(\dpath.RF.R[4][0] ),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(_00074_),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2105 (.A(\dpath.RF.R[22][2] ),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(_00352_),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(\dpath.RF.R[9][20] ),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2108 (.A(_00725_),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(\dpath.RF.R[23][9] ),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\dpath.sd_DX.q[3] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(_00677_),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(\dpath.RF.R[14][2] ),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2112 (.A(_01283_),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(\dpath.RF.R[21][29] ),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(_00443_),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(\dpath.RF.R[31][2] ),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2116 (.A(_00108_),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2117 (.A(\dpath.RF.R[31][24] ),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(_00130_),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(\dpath.RF.R[15][18] ),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_00385_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(_00592_),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(\dpath.RF.R[13][5] ),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2122 (.A(_01478_),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2123 (.A(\dpath.RF.R[15][0] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(_00574_),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(\dpath.RF.R[29][17] ),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(_00155_),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2127 (.A(\dpath.RF.R[27][11] ),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2128 (.A(_00972_),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(\dpath.RF.R[11][23] ),
    .X(net3024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\dpath.RF.R[0][30] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(_00952_),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(\dpath.RF.R[12][8] ),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(_01578_),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2133 (.A(\dpath.RF.R[29][7] ),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(_00145_),
    .X(net3029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(\dpath.RF.R[31][28] ),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(_00134_),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(\dpath.RF.R[15][4] ),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(_00578_),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2139 (.A(\dpath.RF.R[15][10] ),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_00799_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(_00584_),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(\dpath.RF.R[15][1] ),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(_00575_),
    .X(net3037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(\dpath.RF.R[16][26] ),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(_00568_),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2145 (.A(\dpath.RF.R[6][7] ),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(_00049_),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(\dpath.RF.R[31][6] ),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(_00112_),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(\dpath.RF.R[13][10] ),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\dpath.sd_DX.q[5] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(_01483_),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2151 (.A(\dpath.RF.R[7][2] ),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(_00012_),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2153 (.A(\dpath.RF.R[4][23] ),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(_00097_),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(\dpath.RF.R[16][1] ),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(_00543_),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2157 (.A(\dpath.RF.R[24][22] ),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2158 (.A(_01624_),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(\dpath.RF.R[27][25] ),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_00387_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(_00986_),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(\dpath.RF.R[13][0] ),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2162 (.A(_01473_),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(\dpath.RF.R[25][3] ),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(_00740_),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(\dpath.RF.R[21][22] ),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(_00436_),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(\dpath.csrw_out_DX.q[29] ),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(_01470_),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2169 (.A(\dpath.RF.R[13][18] ),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\dpath.RF.R[0][19] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(_01491_),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(\dpath.RF.R[23][23] ),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2172 (.A(_00691_),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2173 (.A(\dpath.RF.R[23][1] ),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(_00669_),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(\dpath.RF.R[4][3] ),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(_00077_),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(\dpath.RF.R[25][11] ),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(_00748_),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2179 (.A(\dpath.RF.R[4][12] ),
    .X(net3074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_00788_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(_00086_),
    .X(net3075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2181 (.A(\dpath.RF.R[31][30] ),
    .X(net3076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(_00136_),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(\dpath.RF.R[29][16] ),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2184 (.A(_00154_),
    .X(net3079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(\dpath.RF.R[31][22] ),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(_00128_),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(\dpath.RF.R[31][3] ),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(_00109_),
    .X(net3083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2189 (.A(\dpath.RF.R[28][0] ),
    .X(net3084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\dpath.RF.R[0][8] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(_00865_),
    .X(net3085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2191 (.A(\ctrl.inst_M[12] ),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(_00303_),
    .X(net3087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(\dpath.RF.R[7][26] ),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(_00036_),
    .X(net3089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(\dpath.RF.R[25][4] ),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(_00741_),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2197 (.A(\dpath.RF.R[11][1] ),
    .X(net3092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(_00930_),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2199 (.A(\dpath.RF.R[25][29] ),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_01193_),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_00777_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(_00766_),
    .X(net3095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(\dpath.RF.R[11][16] ),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2202 (.A(_00945_),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(\dpath.RF.R[20][2] ),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(_00480_),
    .X(net3099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(\dpath.RF.R[21][24] ),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(_00438_),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(\dpath.RF.R[29][12] ),
    .X(net3102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(_00150_),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(\dpath.RF.R[31][5] ),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\ctrl.inst_M[28] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(_00111_),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(\dpath.RF.R[31][26] ),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(_00132_),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(\dpath.RF.R[18][26] ),
    .X(net3108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(_00632_),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2215 (.A(\dpath.RF.R[27][13] ),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(_00974_),
    .X(net3111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(\dpath.RF.R[7][1] ),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(_00011_),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(\dpath.RF.R[11][3] ),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_00314_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(_00932_),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(\ctrl.inst_M[6] ),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(_00297_),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(\dpath.RF.R[3][5] ),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(_00175_),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(\dpath.RF.R[3][20] ),
    .X(net3120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(_00190_),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2227 (.A(\dpath.RF.R[14][1] ),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(_01282_),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(\dpath.RF.R[29][18] ),
    .X(net3124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\dpath.RF.R[0][17] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(_00156_),
    .X(net3125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(\dpath.RF.R[29][14] ),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2232 (.A(_00152_),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(\dpath.RF.R[29][27] ),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(_00165_),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(\dpath.RF.R[7][27] ),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(_00037_),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2237 (.A(\dpath.RF.R[8][30] ),
    .X(net3132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(_01023_),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(\dpath.RF.R[25][5] ),
    .X(net3134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_00786_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(_00742_),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(\dpath.RF.R[23][6] ),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2242 (.A(_00674_),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2243 (.A(\dpath.RF.R[15][20] ),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2244 (.A(_00594_),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2245 (.A(\dpath.RF.R[29][13] ),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(_00151_),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(\dpath.RF.R[27][24] ),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(_00985_),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2249 (.A(\dpath.RF.R[31][27] ),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\dpath.RF.R[0][9] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2250 (.A(_00133_),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(\dpath.RF.R[23][2] ),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2252 (.A(_00670_),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(\dpath.RF.R[27][0] ),
    .X(net3148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2254 (.A(_00961_),
    .X(net3149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(\dpath.RF.R[4][25] ),
    .X(net3150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(_00099_),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(\dpath.RF.R[3][0] ),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(_00170_),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2259 (.A(\dpath.RF.R[23][11] ),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_00778_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(_00679_),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(\dpath.RF.R[13][3] ),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2262 (.A(_01476_),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2263 (.A(\dpath.RF.R[11][11] ),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(_00940_),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2265 (.A(\dpath.RF.R[25][12] ),
    .X(net3160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(_00749_),
    .X(net3161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2267 (.A(\dpath.RF.R[27][19] ),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(_00980_),
    .X(net3163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(\dpath.RF.R[11][30] ),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\dpath.RF.R[0][31] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(_00959_),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2271 (.A(\dpath.RF.R[5][26] ),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(_00228_),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(\dpath.RF.R[31][11] ),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2274 (.A(_00117_),
    .X(net3169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(\dpath.csrw_out_DX.q[2] ),
    .X(net3170));
 sky130_fd_sc_hd__buf_1 hold2276 (.A(_01443_),
    .X(net3171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(\dpath.RF.R[29][11] ),
    .X(net3172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2278 (.A(_00149_),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2279 (.A(\dpath.RF.R[31][25] ),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_00800_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(_00131_),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2281 (.A(\ctrl.d2c_inst[3] ),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(_00267_),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2283 (.A(\dpath.csrw_out_DX.q[7] ),
    .X(net3178));
 sky130_fd_sc_hd__buf_1 hold2284 (.A(_01448_),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2285 (.A(\dpath.RF.R[29][0] ),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(_00138_),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(\dpath.RF.R[31][8] ),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(_00114_),
    .X(net3183));
 sky130_fd_sc_hd__buf_1 hold2289 (.A(net3726),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\dpath.RF.R[0][10] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(_01440_),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(\dpath.RF.R[3][6] ),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(_00176_),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(\dpath.RF.R[22][6] ),
    .X(net3188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(_00356_),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(\dpath.RF.R[13][13] ),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(_01486_),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(\dpath.RF.R[4][26] ),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(_00100_),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2299 (.A(\dpath.csrw_out_DX.q[3] ),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\dpath.csrw_out_DX.q[25] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_00779_),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_2 hold2300 (.A(_01444_),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2301 (.A(\dpath.RF.R[23][26] ),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(_00694_),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(\ctrl.val_M ),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(_00235_),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(\ctrl.inst_M[10] ),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2306 (.A(_01783_),
    .X(net3201));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2307 (.A(net3736),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(\ctrl.inst_M[8] ),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(_01781_),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\dpath.RF.R[0][14] ),
    .X(net1126));
 sky130_fd_sc_hd__buf_1 hold2310 (.A(net3725),
    .X(net3205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(\dpath.sd_DX.q[10] ),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2312 (.A(\ctrl.inst_X[4] ),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2313 (.A(\ctrl.inst_M[2] ),
    .X(net3208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(\ctrl.inst_X[5] ),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2315 (.A(\dpath.csrw_out_DX.q[6] ),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(\ctrl.d2c_inst[2] ),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(\ctrl.inst_M[3] ),
    .X(net3212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2318 (.A(_00294_),
    .X(net3213));
 sky130_fd_sc_hd__clkbuf_2 hold2319 (.A(\dpath.csrw_out0.d[0] ),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_00783_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(_01089_),
    .X(net3215));
 sky130_fd_sc_hd__clkbuf_2 hold2321 (.A(net3751),
    .X(net3216));
 sky130_fd_sc_hd__buf_2 hold2322 (.A(\dpath.csrw_out0.d[24] ),
    .X(net3217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(_01113_),
    .X(net3218));
 sky130_fd_sc_hd__buf_1 hold2324 (.A(net3728),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(\dpath.csrw_out_DX.q[9] ),
    .X(net3220));
 sky130_fd_sc_hd__buf_1 hold2326 (.A(\dpath.inst_pc[17] ),
    .X(net3221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(_01523_),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(\dpath.btarg_DX.q[30] ),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(_05676_),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\dpath.sd_DX.q[4] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(_00666_),
    .X(net3225));
 sky130_fd_sc_hd__buf_1 hold2331 (.A(\ctrl.d2c_inst[16] ),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(_01635_),
    .X(net3227));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2333 (.A(net3752),
    .X(net3228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(_01418_),
    .X(net3229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(\dpath.csrw_out_DX.q[4] ),
    .X(net3230));
 sky130_fd_sc_hd__buf_1 hold2336 (.A(net3742),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(_01509_),
    .X(net3232));
 sky130_fd_sc_hd__buf_1 hold2338 (.A(net3763),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(_01507_),
    .X(net3234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_00386_),
    .X(net1129));
 sky130_fd_sc_hd__buf_1 hold2340 (.A(net3727),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(\ctrl.inst_M[5] ),
    .X(net3236));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2342 (.A(net3741),
    .X(net3237));
 sky130_fd_sc_hd__buf_1 hold2343 (.A(net3745),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2344 (.A(_01510_),
    .X(net3239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2345 (.A(\ctrl.inst_M[7] ),
    .X(net3240));
 sky130_fd_sc_hd__buf_1 hold2346 (.A(\dpath.inst_pc[15] ),
    .X(net3241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2347 (.A(_01521_),
    .X(net3242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(\ctrl.inst_X[8] ),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(\dpath.sd_DX.q[29] ),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\dpath.RF.R[0][13] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(\ctrl.inst_X[9] ),
    .X(net3245));
 sky130_fd_sc_hd__buf_1 hold2351 (.A(net3756),
    .X(net3246));
 sky130_fd_sc_hd__buf_2 hold2352 (.A(\dpath.csrw_out0.d[18] ),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(_01107_),
    .X(net3248));
 sky130_fd_sc_hd__buf_1 hold2354 (.A(net3739),
    .X(net3249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2355 (.A(_06880_),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(_06881_),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(\dpath.btarg_DX.q[27] ),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(_05118_),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(_00663_),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_00782_),
    .X(net1131));
 sky130_fd_sc_hd__buf_2 hold2360 (.A(\dpath.csrw_out0.d[23] ),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(_01112_),
    .X(net3256));
 sky130_fd_sc_hd__clkbuf_2 hold2362 (.A(\dpath.csrw_out0.d[1] ),
    .X(net3257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2363 (.A(_01090_),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2364 (.A(\ctrl.inst_M[4] ),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(\dpath.btarg_DX.q[0] ),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(_01746_),
    .X(net3261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(_01671_),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(\ctrl.d2c_inst[5] ),
    .X(net3263));
 sky130_fd_sc_hd__buf_1 hold2369 (.A(net3738),
    .X(net3264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\ctrl.inst_M[13] ),
    .X(net1132));
 sky130_fd_sc_hd__buf_1 hold2370 (.A(net3754),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2371 (.A(_01522_),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2372 (.A(\dpath.RF.wdata[4] ),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(_02218_),
    .X(net3268));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2374 (.A(_02247_),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2375 (.A(\dpath.sd_DX.q[30] ),
    .X(net3270));
 sky130_fd_sc_hd__buf_1 hold2376 (.A(\dpath.RF.wdata[3] ),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(_02164_),
    .X(net3272));
 sky130_fd_sc_hd__clkbuf_2 hold2378 (.A(_02184_),
    .X(net3273));
 sky130_fd_sc_hd__buf_1 hold2379 (.A(net3750),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_00304_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(_01516_),
    .X(net3275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2381 (.A(\ctrl.d2c_inst[2] ),
    .X(net3276));
 sky130_fd_sc_hd__buf_1 hold2382 (.A(net3735),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2383 (.A(_01513_),
    .X(net3278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(\ctrl.inst_X[11] ),
    .X(net3279));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2385 (.A(net255),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(\ctrl.inst_X[10] ),
    .X(net3281));
 sky130_fd_sc_hd__buf_1 hold2387 (.A(net3737),
    .X(net3282));
 sky130_fd_sc_hd__buf_1 hold2388 (.A(\dpath.inst_pc[30] ),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(_01536_),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\dpath.RF.R[0][18] ),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_2 hold2390 (.A(net3746),
    .X(net3285));
 sky130_fd_sc_hd__buf_1 hold2391 (.A(net3744),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(_01514_),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2393 (.A(\dpath.sd_DX.q[26] ),
    .X(net3288));
 sky130_fd_sc_hd__clkbuf_2 hold2394 (.A(\dpath.csrw_out0.d[31] ),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(_01120_),
    .X(net3290));
 sky130_fd_sc_hd__buf_1 hold2396 (.A(net3748),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(_01520_),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(net298),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(_01072_),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_01466_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_00787_),
    .X(net1135));
 sky130_fd_sc_hd__buf_1 hold2400 (.A(\dpath.inst_pc[13] ),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2401 (.A(_01519_),
    .X(net3296));
 sky130_fd_sc_hd__buf_1 hold2402 (.A(net3740),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2403 (.A(_01512_),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(net299),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(_01073_),
    .X(net3300));
 sky130_fd_sc_hd__buf_1 hold2406 (.A(net3734),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2407 (.A(_01518_),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(net301),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(_01075_),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\dpath.RF.R[0][26] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(net333),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2411 (.A(_05879_),
    .X(net3306));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2412 (.A(\ctrl.inst_X[21] ),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(\dpath.sd_DX.q[31] ),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(\ctrl.inst_X[7] ),
    .X(net3309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(\dpath.RF.wdata[0] ),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2416 (.A(_05991_),
    .X(net3311));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2417 (.A(\ctrl.inst_X[23] ),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2418 (.A(net297),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(_01071_),
    .X(net3314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_00795_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2420 (.A(net296),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(_01070_),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(net295),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(_01069_),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2424 (.A(net294),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2425 (.A(_01068_),
    .X(net3320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2426 (.A(net302),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(_01076_),
    .X(net3322));
 sky130_fd_sc_hd__buf_1 hold2428 (.A(\dpath.inst_pc[19] ),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(_01525_),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\ctrl.inst_M[29] ),
    .X(net1138));
 sky130_fd_sc_hd__buf_1 hold2430 (.A(\dpath.inst_pc[18] ),
    .X(net3325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2431 (.A(_01524_),
    .X(net3326));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2432 (.A(\ctrl.val_DX.q ),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(net320),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(_01063_),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(net322),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(_01065_),
    .X(net3331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(net300),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(_01074_),
    .X(net3333));
 sky130_fd_sc_hd__clkbuf_2 hold2439 (.A(\dpath.csrw_out0.d[17] ),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_00315_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(_01106_),
    .X(net3335));
 sky130_fd_sc_hd__buf_1 hold2441 (.A(\dpath.csrr[30] ),
    .X(net3336));
 sky130_fd_sc_hd__clkbuf_2 hold2442 (.A(_05662_),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(_01439_),
    .X(net3338));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2444 (.A(net3755),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(_01436_),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(net228),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(\ctrl.d2c_inst[14] ),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(net321),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(_01064_),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\dpath.csrw_out_DX.q[0] ),
    .X(net1140));
 sky130_fd_sc_hd__buf_1 hold2450 (.A(net3743),
    .X(net3345));
 sky130_fd_sc_hd__buf_1 hold2451 (.A(\dpath.csrr[12] ),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(net318),
    .X(net3347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(_01061_),
    .X(net3348));
 sky130_fd_sc_hd__clkbuf_2 hold2454 (.A(net3753),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2455 (.A(net305),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(_01078_),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(net293),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2458 (.A(_01067_),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(net308),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_01441_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(_01081_),
    .X(net3355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(net309),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2462 (.A(_01082_),
    .X(net3357));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2463 (.A(net3747),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2464 (.A(_01420_),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(net306),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(_01079_),
    .X(net3361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(net307),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2468 (.A(_01080_),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2469 (.A(net323),
    .X(net3364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\dpath.RF.R[0][12] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(_01066_),
    .X(net3365));
 sky130_fd_sc_hd__clkbuf_2 hold2471 (.A(\dpath.csrw_out0.d[16] ),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2472 (.A(_01105_),
    .X(net3367));
 sky130_fd_sc_hd__buf_1 hold2473 (.A(net246),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(_00662_),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2475 (.A(net304),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2476 (.A(_01077_),
    .X(net3371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(\dpath.btarg_DX.q[21] ),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(_04122_),
    .X(net3373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2479 (.A(_00657_),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_00781_),
    .X(net1143));
 sky130_fd_sc_hd__buf_1 hold2480 (.A(net259),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(net314),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(_01059_),
    .X(net3377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(net315),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2484 (.A(_01087_),
    .X(net3379));
 sky130_fd_sc_hd__buf_2 hold2485 (.A(\dpath.csrw_out0.d[27] ),
    .X(net3380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(_01116_),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2487 (.A(net292),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(_01057_),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(net312),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\dpath.RF.R[0][15] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2490 (.A(_01085_),
    .X(net3385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(net311),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2492 (.A(_01084_),
    .X(net3387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(net310),
    .X(net3388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2494 (.A(_01083_),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(net319),
    .X(net3390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(_01062_),
    .X(net3391));
 sky130_fd_sc_hd__clkbuf_4 hold2497 (.A(\ctrl.d2c_inst[25] ),
    .X(net3392));
 sky130_fd_sc_hd__clkbuf_2 hold2498 (.A(\ctrl.d2c_inst[21] ),
    .X(net3393));
 sky130_fd_sc_hd__buf_1 hold2499 (.A(net244),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\dpath.csrw_out_MW.d[16] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_00784_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2500 (.A(_00660_),
    .X(net3395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2501 (.A(\dpath.btarg_DX.q[22] ),
    .X(net3396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2502 (.A(_04280_),
    .X(net3397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(_00658_),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2504 (.A(\dpath.csrr[7] ),
    .X(net3399));
 sky130_fd_sc_hd__clkbuf_2 hold2505 (.A(_02460_),
    .X(net3400));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2506 (.A(\dpath.inst_pc[28] ),
    .X(net3401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(_01534_),
    .X(net3402));
 sky130_fd_sc_hd__clkbuf_2 hold2508 (.A(net3758),
    .X(net3403));
 sky130_fd_sc_hd__clkbuf_2 hold2509 (.A(\dpath.csrw_out0.d[15] ),
    .X(net3404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\dpath.RF.R[0][1] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2510 (.A(_01104_),
    .X(net3405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(net303),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(_01058_),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(net317),
    .X(net3408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2514 (.A(_01060_),
    .X(net3409));
 sky130_fd_sc_hd__buf_1 hold2515 (.A(net230),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2516 (.A(net190),
    .X(net3411));
 sky130_fd_sc_hd__buf_1 hold2517 (.A(_02388_),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(net313),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2519 (.A(_01086_),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_00770_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(_02009_),
    .X(net3415));
 sky130_fd_sc_hd__buf_1 hold2521 (.A(\dpath.csrr[8] ),
    .X(net3416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(_02552_),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2523 (.A(net316),
    .X(net3418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(_01088_),
    .X(net3419));
 sky130_fd_sc_hd__clkbuf_4 hold2525 (.A(\ctrl.d2c_inst[27] ),
    .X(net3420));
 sky130_fd_sc_hd__clkbuf_4 hold2526 (.A(\ctrl.d2c_inst[28] ),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(\dpath.btarg_DX.q[31] ),
    .X(net3422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2528 (.A(_05836_),
    .X(net3423));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2529 (.A(\ctrl.inst_X[22] ),
    .X(net3424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\dpath.RF.R[0][11] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2530 (.A(\dpath.sd_DX.q[27] ),
    .X(net3425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(\dpath.btarg_DX.q[11] ),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(_02851_),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(_02852_),
    .X(net3428));
 sky130_fd_sc_hd__buf_1 hold2534 (.A(net3749),
    .X(net3429));
 sky130_fd_sc_hd__buf_2 hold2535 (.A(\dpath.csrw_out0.d[26] ),
    .X(net3430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(_01115_),
    .X(net3431));
 sky130_fd_sc_hd__clkbuf_2 hold2537 (.A(\ctrl.d2c_inst[20] ),
    .X(net3432));
 sky130_fd_sc_hd__clkbuf_2 hold2538 (.A(\dpath.csrw_out0.d[13] ),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(_01102_),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_00780_),
    .X(net1149));
 sky130_fd_sc_hd__clkbuf_4 hold2540 (.A(\ctrl.d2c_inst[30] ),
    .X(net3435));
 sky130_fd_sc_hd__clkbuf_2 hold2541 (.A(net3761),
    .X(net3436));
 sky130_fd_sc_hd__buf_2 hold2542 (.A(\dpath.csrw_out0.d[29] ),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(_01118_),
    .X(net3438));
 sky130_fd_sc_hd__clkbuf_2 hold2544 (.A(net3730),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(_01438_),
    .X(net3440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2546 (.A(net247),
    .X(net3441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(\dpath.sd_DX.q[28] ),
    .X(net3442));
 sky130_fd_sc_hd__clkbuf_2 hold2548 (.A(\dpath.csrw_out0.d[2] ),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(_01091_),
    .X(net3444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\ctrl.inst_X[3] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2550 (.A(net331),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2551 (.A(_05877_),
    .X(net3446));
 sky130_fd_sc_hd__buf_1 hold2552 (.A(net249),
    .X(net3447));
 sky130_fd_sc_hd__buf_2 hold2553 (.A(\dpath.csrw_out0.d[22] ),
    .X(net3448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(_01111_),
    .X(net3449));
 sky130_fd_sc_hd__buf_2 hold2555 (.A(\dpath.csrw_out0.d[25] ),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(_01114_),
    .X(net3451));
 sky130_fd_sc_hd__buf_2 hold2557 (.A(\ctrl.d2c_inst[26] ),
    .X(net3452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(\dpath.csrr[16] ),
    .X(net3453));
 sky130_fd_sc_hd__clkbuf_2 hold2559 (.A(_03412_),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_00239_),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_2 hold2560 (.A(net3757),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2561 (.A(_01527_),
    .X(net3456));
 sky130_fd_sc_hd__buf_2 hold2562 (.A(\dpath.csrw_out0.d[14] ),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(_01103_),
    .X(net3458));
 sky130_fd_sc_hd__buf_2 hold2564 (.A(\dpath.csrw_out0.d[28] ),
    .X(net3459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2565 (.A(_01117_),
    .X(net3460));
 sky130_fd_sc_hd__clkbuf_4 hold2566 (.A(\ctrl.d2c_inst[29] ),
    .X(net3461));
 sky130_fd_sc_hd__clkbuf_2 hold2567 (.A(\dpath.inst_pc[20] ),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2568 (.A(_01526_),
    .X(net3463));
 sky130_fd_sc_hd__buf_1 hold2569 (.A(net3760),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\ctrl.inst_M[27] ),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_2 hold2570 (.A(net3759),
    .X(net3465));
 sky130_fd_sc_hd__clkbuf_2 hold2571 (.A(\dpath.inst_pc[22] ),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2572 (.A(_01528_),
    .X(net3467));
 sky130_fd_sc_hd__clkbuf_2 hold2573 (.A(\dpath.inst_pc[23] ),
    .X(net3468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(_01529_),
    .X(net3469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(\ctrl.d2c_inst[12] ),
    .X(net3470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2576 (.A(net248),
    .X(net3471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2577 (.A(_00664_),
    .X(net3472));
 sky130_fd_sc_hd__buf_1 hold2578 (.A(net258),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(_00644_),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_00313_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(\dpath.btarg_DX.q[2] ),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(_02141_),
    .X(net3476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2582 (.A(_00638_),
    .X(net3477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(\dpath.btarg_DX.q[4] ),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(_02259_),
    .X(net3479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2585 (.A(_00640_),
    .X(net3480));
 sky130_fd_sc_hd__buf_2 hold2586 (.A(\dpath.csrw_out0.d[3] ),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(_01092_),
    .X(net3482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2588 (.A(\dpath.csrr[10] ),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(_02734_),
    .X(net3484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\dpath.RF.R[0][28] ),
    .X(net1154));
 sky130_fd_sc_hd__buf_1 hold2590 (.A(_02741_),
    .X(net3485));
 sky130_fd_sc_hd__buf_2 hold2591 (.A(\dpath.csrw_out0.d[20] ),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(_01109_),
    .X(net3487));
 sky130_fd_sc_hd__buf_2 hold2593 (.A(\dpath.csrw_out0.d[19] ),
    .X(net3488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(_01108_),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(\ctrl.d2c_inst[20] ),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(\dpath.btarg_DX.q[29] ),
    .X(net3491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2597 (.A(_00665_),
    .X(net3492));
 sky130_fd_sc_hd__buf_1 hold2598 (.A(net253),
    .X(net3493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(_00639_),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_01201_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_00797_),
    .X(net1155));
 sky130_fd_sc_hd__buf_1 hold2600 (.A(net3762),
    .X(net3495));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2601 (.A(\ctrl.d2c_inst[17] ),
    .X(net3496));
 sky130_fd_sc_hd__buf_2 hold2602 (.A(\dpath.csrw_out0.d[8] ),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(_01097_),
    .X(net3498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(\ctrl.d2c_inst[5] ),
    .X(net3499));
 sky130_fd_sc_hd__buf_2 hold2605 (.A(\dpath.csrw_out0.d[21] ),
    .X(net3500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(_01110_),
    .X(net3501));
 sky130_fd_sc_hd__buf_2 hold2607 (.A(\dpath.csrw_out0.d[9] ),
    .X(net3502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(_01098_),
    .X(net3503));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2609 (.A(\dpath.csrr[14] ),
    .X(net3504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\ctrl.inst_X[12] ),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_2 hold2610 (.A(\dpath.csrw_out0.d[30] ),
    .X(net3505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2611 (.A(_01119_),
    .X(net3506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(net245),
    .X(net3507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(_00661_),
    .X(net3508));
 sky130_fd_sc_hd__clkbuf_2 hold2614 (.A(net3729),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(net234),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(_00651_),
    .X(net3511));
 sky130_fd_sc_hd__buf_2 hold2617 (.A(\dpath.csrw_out0.d[10] ),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(_01099_),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(net257),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_01763_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(_00643_),
    .X(net3515));
 sky130_fd_sc_hd__buf_2 hold2621 (.A(\dpath.csrw_out0.d[5] ),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(_01094_),
    .X(net3517));
 sky130_fd_sc_hd__buf_1 hold2623 (.A(\dpath.inst_pc[2] ),
    .X(net3518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2624 (.A(_01688_),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(net262),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2626 (.A(_01100_),
    .X(net3521));
 sky130_fd_sc_hd__clkbuf_2 hold2627 (.A(net3731),
    .X(net3522));
 sky130_fd_sc_hd__buf_2 hold2628 (.A(\dpath.csrw_out0.d[4] ),
    .X(net3523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(_01093_),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\dpath.RF.R[0][5] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(net238),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(_00655_),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2632 (.A(net239),
    .X(net3527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(_01672_),
    .X(net3528));
 sky130_fd_sc_hd__buf_2 hold2634 (.A(\dpath.csrw_out0.d[7] ),
    .X(net3529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(_01096_),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2636 (.A(\ctrl.d2c_inst[3] ),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2637 (.A(net263),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2638 (.A(_01101_),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(\dpath.btarg_DX.q[5] ),
    .X(net3534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_00774_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(_02325_),
    .X(net3535));
 sky130_fd_sc_hd__buf_1 hold2641 (.A(\ctrl.d2c_inst[18] ),
    .X(net3536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2642 (.A(net240),
    .X(net3537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(_00656_),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(net232),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(_00649_),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2646 (.A(net173),
    .X(net3541));
 sky130_fd_sc_hd__clkbuf_2 hold2647 (.A(net3732),
    .X(net3542));
 sky130_fd_sc_hd__buf_1 hold2648 (.A(\dpath.csrr[4] ),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(net236),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\dpath.RF.R[0][29] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2650 (.A(_00653_),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(net243),
    .X(net3546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(_00659_),
    .X(net3547));
 sky130_fd_sc_hd__buf_2 hold2653 (.A(\dpath.csrw_out0.d[6] ),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(_01095_),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(\ctrl.d2c_inst[4] ),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(net326),
    .X(net3551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(_05872_),
    .X(net3552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(net354),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2659 (.A(net353),
    .X(net3554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_00798_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2660 (.A(net233),
    .X(net3555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(_00650_),
    .X(net3556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2662 (.A(net351),
    .X(net3557));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2663 (.A(net235),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(_00652_),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2665 (.A(net335),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(_05862_),
    .X(net3561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(net352),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(net349),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(_05864_),
    .X(net3564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\ctrl.inst_M[30] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(\dpath.btarg_DX.q[9] ),
    .X(net3565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(net350),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(net327),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(_05873_),
    .X(net3568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(net330),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(_05876_),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(net324),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(_05861_),
    .X(net3572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(net332),
    .X(net3573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(_05878_),
    .X(net3574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_00316_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(net237),
    .X(net3575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(_00654_),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2682 (.A(net325),
    .X(net3577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(_05871_),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(net231),
    .X(net3579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2685 (.A(_00648_),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(net355),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(\dpath.btarg_DX.q[6] ),
    .X(net3582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(_02396_),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2689 (.A(_00642_),
    .X(net3584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\dpath.RF.R[0][23] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2690 (.A(net336),
    .X(net3585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(\dpath.RF.wdata[13] ),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2692 (.A(net229),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2693 (.A(_00646_),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2694 (.A(net184),
    .X(net3589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(net179),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(net348),
    .X(net3591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2697 (.A(_05892_),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2698 (.A(net339),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(net343),
    .X(net3594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\ctrl.inst_M[23] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_00792_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(net337),
    .X(net3595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(net347),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(_05891_),
    .X(net3597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(net171),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(net340),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(net338),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(\dpath.csrr[26] ),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(_04933_),
    .X(net3602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(net346),
    .X(net3603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2709 (.A(_05863_),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\ctrl.inst_X[2] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2710 (.A(net162),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2711 (.A(net172),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(net334),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2713 (.A(net345),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(\dpath.csrr[28] ),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(_05292_),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2716 (.A(net342),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2717 (.A(_05887_),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2718 (.A(net329),
    .X(net3613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(_05875_),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_00238_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(net341),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(_05886_),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2722 (.A(net344),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(_05889_),
    .X(net3618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(net328),
    .X(net3619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2725 (.A(_05874_),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2726 (.A(net166),
    .X(net3621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(net176),
    .X(net3622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(\dpath.RF.wdata[21] ),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(net189),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\ctrl.inst_M[14] ),
    .X(net1168));
 sky130_fd_sc_hd__buf_1 hold2730 (.A(_06182_),
    .X(net3625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(\dpath.csrr[23] ),
    .X(net3626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2732 (.A(\dpath.RF.wdata[11] ),
    .X(net3627));
 sky130_fd_sc_hd__buf_1 hold2733 (.A(_02775_),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2734 (.A(_02841_),
    .X(net3629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(\dpath.RF.wdata[20] ),
    .X(net3630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(\dpath.csrr[22] ),
    .X(net3631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(net178),
    .X(net3632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2738 (.A(net170),
    .X(net3633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(net168),
    .X(net3634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_00305_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2740 (.A(\dpath.alu.adder.in1[26] ),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2741 (.A(net177),
    .X(net3636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(\dpath.RF.wdata[28] ),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(net165),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(net167),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(net193),
    .X(net3640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(net163),
    .X(net3641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(net169),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(net174),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2749 (.A(\dpath.RF.wdata[24] ),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\dpath.RF.R[0][2] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2750 (.A(net192),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(\dpath.csrr[27] ),
    .X(net3646));
 sky130_fd_sc_hd__buf_1 hold2752 (.A(_05109_),
    .X(net3647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(net164),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(\dpath.csrr[19] ),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2755 (.A(net187),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(net188),
    .X(net3651));
 sky130_fd_sc_hd__buf_1 hold2757 (.A(\dpath.csrr[0] ),
    .X(net3652));
 sky130_fd_sc_hd__buf_1 hold2758 (.A(\dpath.csrr[5] ),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(net191),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_00771_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2760 (.A(net180),
    .X(net3655));
 sky130_fd_sc_hd__buf_1 hold2761 (.A(\dpath.csrr[6] ),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(\dpath.csrr[15] ),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(net175),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(\dpath.RF.wdata[26] ),
    .X(net3659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(net665),
    .X(net3660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(_06687_),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(\dpath.csrr[9] ),
    .X(net3662));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2768 (.A(net183),
    .X(net3663));
 sky130_fd_sc_hd__buf_1 hold2769 (.A(net186),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\ctrl.inst_M[9] ),
    .X(net1172));
 sky130_fd_sc_hd__clkbuf_4 hold2770 (.A(_00004_),
    .X(net3665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(_06780_),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(net181),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(\dpath.csrr[20] ),
    .X(net3668));
 sky130_fd_sc_hd__clkbuf_2 hold2774 (.A(_00003_),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(_06725_),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(_06732_),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(\dpath.csrr[17] ),
    .X(net3672));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2778 (.A(_03543_),
    .X(net3673));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2779 (.A(\dpath.csrr[29] ),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_01782_),
    .X(net1173));
 sky130_fd_sc_hd__clkbuf_2 hold2780 (.A(_05476_),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(net182),
    .X(net3676));
 sky130_fd_sc_hd__buf_1 hold2782 (.A(_00004_),
    .X(net3677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(\dpath.RF.wdata[5] ),
    .X(net3678));
 sky130_fd_sc_hd__buf_1 hold2784 (.A(\dpath.csrr[31] ),
    .X(net3679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(_05828_),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(net185),
    .X(net3681));
 sky130_fd_sc_hd__buf_1 hold2787 (.A(\dpath.csrr[1] ),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2788 (.A(\dpath.csrr[3] ),
    .X(net3683));
 sky130_fd_sc_hd__buf_1 hold2789 (.A(\dpath.csrr[2] ),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\dpath.RF.R[0][24] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2790 (.A(\dpath.csrr[11] ),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(\dpath.csrr[21] ),
    .X(net3686));
 sky130_fd_sc_hd__buf_1 hold2792 (.A(\dpath.csrr[24] ),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(\dpath.csrr[13] ),
    .X(net3688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(\dpath.RF.wdata[29] ),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(\dpath.csrr[18] ),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(\dpath.csrr[25] ),
    .X(net3691));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2797 (.A(_04759_),
    .X(net3692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(\dpath.RF.R[21][14] ),
    .X(net3693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2799 (.A(\dpath.RF.R[27][10] ),
    .X(net3694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_00309_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_00793_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2800 (.A(\dpath.RF.R[24][24] ),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(\dpath.RF.wdata[14] ),
    .X(net3696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(\dpath.RF.R[21][6] ),
    .X(net3697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2803 (.A(\dpath.RF.R[31][1] ),
    .X(net3698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(_06071_),
    .X(net3699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(\dpath.RF.R[22][17] ),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(_06455_),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(_06460_),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2808 (.A(\dpath.RF.R[22][9] ),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2809 (.A(\dpath.RF.wdata[28] ),
    .X(net3704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\ctrl.inst_X[0] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2810 (.A(\dpath.RF.R[20][16] ),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(\dpath.RF.R[26][21] ),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2812 (.A(_06545_),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2813 (.A(\dpath.RF.R[25][2] ),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2814 (.A(\dpath.RF.R[19][8] ),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(\dpath.RF.R[28][6] ),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(\dpath.RF.wdata[1] ),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(\dpath.RF.wdata[30] ),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(\dpath.RF.R[21][19] ),
    .X(net3713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2819 (.A(\dpath.RF.wdata[22] ),
    .X(net3714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_00236_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2820 (.A(\ctrl.d2c_inst[14] ),
    .X(net3715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2821 (.A(\dpath.RF.wdata[14] ),
    .X(net3716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(\dpath.RF.wdata[12] ),
    .X(net3717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(\dpath.RF.wdata[14] ),
    .X(net3718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(\ctrl.d2c_inst[7] ),
    .X(net3725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(\dpath.inst_pc[31] ),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(\ctrl.d2c_inst[8] ),
    .X(net3727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(\ctrl.d2c_inst[11] ),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(\dpath.inst_pc[26] ),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(\dpath.inst_pc[29] ),
    .X(net3730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\dpath.RF.R[0][16] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(\dpath.inst_pc[25] ),
    .X(net3731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(\dpath.inst_pc[24] ),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2832 (.A(\dpath.inst_pc[5] ),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(\dpath.inst_pc[12] ),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(\dpath.inst_pc[7] ),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2835 (.A(\ctrl.d2c_inst[9] ),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(\ctrl.d2c_inst[13] ),
    .X(net3737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(\ctrl.d2c_inst[12] ),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2838 (.A(\dpath.inst_pc[0] ),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(\dpath.inst_pc[6] ),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_00785_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2840 (.A(\ctrl.d2c_inst[10] ),
    .X(net3741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(\dpath.inst_pc[3] ),
    .X(net3742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(\ctrl.d2c_inst[6] ),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(\dpath.inst_pc[8] ),
    .X(net3744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(\dpath.inst_pc[4] ),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2845 (.A(\ctrl.d2c_inst[23] ),
    .X(net3746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2846 (.A(\dpath.inst_pc[11] ),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2847 (.A(\dpath.inst_pc[14] ),
    .X(net3748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(\ctrl.d2c_inst[4] ),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(\dpath.inst_pc[10] ),
    .X(net3750));
 sky130_fd_sc_hd__buf_1 hold285 (.A(\dpath.RF.wdata[8] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(\ctrl.d2c_inst[31] ),
    .X(net3751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(\dpath.inst_pc[9] ),
    .X(net3752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(\ctrl.d2c_inst[24] ),
    .X(net3753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(\dpath.inst_pc[16] ),
    .X(net3754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2854 (.A(\dpath.inst_pc[27] ),
    .X(net3755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(net252),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(\dpath.inst_pc[21] ),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2857 (.A(\ctrl.d2c_inst[22] ),
    .X(net3758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(\ctrl.val_D ),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2859 (.A(\ctrl.d2c_inst[15] ),
    .X(net3760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_00326_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(\ctrl.inst_X[20] ),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2861 (.A(\ctrl.d2c_inst[19] ),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2862 (.A(\dpath.inst_pc[1] ),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\dpath.RF.R[8][29] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_01022_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\dpath.RF.R[9][0] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ctrl.inst_M[21] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_00705_),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\dpath.RF.R[5][17] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_00219_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\dpath.RF.R[5][28] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_00230_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\dpath.RF.R[10][25] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_00858_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\dpath.RF.R[1][24] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_00534_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\dpath.RF.R[8][25] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\dpath.csrw_out_DX.q[12] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00307_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_01018_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\dpath.RF.R[1][2] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_00512_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\dpath.RF.R[5][12] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_00214_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\dpath.RF.R[22][18] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_00368_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\dpath.RF.R[14][20] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_01301_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\dpath.RF.R[18][27] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\dpath.csrw_out_MW.d[9] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_00633_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\dpath.RF.R[2][24] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_00825_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\ctrl.inst_X[1] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_00237_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\dpath.RF.R[12][26] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_01596_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\dpath.RF.R[1][28] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_00538_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\dpath.RF.R[16][10] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_01194_),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_00552_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\ctrl.inst_M[26] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_00312_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\dpath.RF.R[10][21] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_00854_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\dpath.RF.R[26][23] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_00920_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\dpath.RF.R[17][2] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_00448_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\dpath.RF.R[30][23] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\dpath.csrw_out_MW.d[22] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_01662_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\dpath.RF.R[26][25] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_00922_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\dpath.RF.R[1][6] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_00516_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\dpath.RF.R[1][23] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_00533_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\dpath.RF.R[16][6] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_00548_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\dpath.RF.R[12][9] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_01207_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_01579_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\dpath.RF.R[10][30] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_00863_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\dpath.RF.R[26][1] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_00898_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\dpath.RF.R[1][7] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_00517_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\dpath.RF.R[14][17] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_01298_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\dpath.RF.R[9][28] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\dpath.csrw_out_DX.q[19] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_00733_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\dpath.RF.R[10][17] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_00850_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\dpath.RF.R[2][30] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_00831_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\dpath.RF.R[30][24] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_01663_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\dpath.RF.R[22][30] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_00380_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\dpath.RF.R[22][3] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_01460_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_00353_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\dpath.RF.R[30][31] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_01670_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\dpath.RF.R[10][28] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_00861_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\dpath.RF.R[1][12] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_00522_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\dpath.RF.R[12][31] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_01601_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\dpath.RF.R[8][31] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\ctrl.inst_M[22] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_01024_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\dpath.RF.R[8][28] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_01021_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\dpath.RF.R[12][17] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_01587_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\dpath.RF.R[10][8] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_00841_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\dpath.RF.R[12][20] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_01590_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\dpath.RF.R[20][8] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_00308_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_00486_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\dpath.RF.R[18][3] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_00609_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\dpath.RF.R[16][21] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_00563_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\dpath.RF.R[9][31] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_00736_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\dpath.RF.R[5][5] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_00207_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\dpath.RF.R[22][21] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\dpath.csrw_out_MW.d[19] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_00371_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\dpath.RF.R[22][0] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_00350_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\dpath.RF.R[14][25] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_01306_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\dpath.RF.R[30][16] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_01655_),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\dpath.RF.R[6][21] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_00063_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\dpath.RF.R[30][30] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_01453_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_01204_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_01669_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\dpath.RF.R[5][30] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_00232_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\dpath.RF.R[1][3] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_00513_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\dpath.RF.R[24][16] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_01618_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\dpath.RF.R[16][20] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_00562_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\dpath.RF.R[18][8] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\dpath.csrw_out_DX.q[24] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_00614_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\dpath.RF.R[14][28] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_01309_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\dpath.RF.R[9][29] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_00734_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\dpath.RF.R[16][5] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_00547_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\dpath.RF.R[22][19] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_00369_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\dpath.RF.R[24][25] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_01465_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_01627_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\dpath.RF.R[5][8] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_00210_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\dpath.RF.R[20][3] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_00481_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\dpath.RF.R[20][24] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_00502_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\dpath.RF.R[30][18] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_01657_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\dpath.RF.R[26][10] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\dpath.csrw_out_DX.q[28] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_00907_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\dpath.RF.R[9][25] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_00730_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\dpath.RF.R[17][26] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_00472_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\dpath.RF.R[28][5] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_00870_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\dpath.RF.R[30][25] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_01664_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\dpath.RF.R[25][0] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_01469_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_00737_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\dpath.RF.R[18][7] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_00613_),
    .X(net1337));
 sky130_fd_sc_hd__buf_1 hold443 (.A(net3733),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_01414_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\dpath.RF.R[28][22] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_00887_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\dpath.RF.R[12][21] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_01591_),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\dpath.RF.R[13][26] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\dpath.csrw_out_MW.d[5] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_01499_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\dpath.RF.R[14][30] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_01311_),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\dpath.RF.R[28][2] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_00867_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\dpath.RF.R[8][19] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_01012_),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\dpath.RF.R[15][8] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_00582_),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\dpath.RF.R[12][13] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_01190_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_01583_),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\dpath.RF.R[16][8] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_00550_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\dpath.RF.R[16][15] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_00557_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\dpath.RF.wdata[6] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_00871_),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\dpath.RF.R[22][24] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_00374_),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\dpath.RF.R[28][31] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\dpath.csrw_out_MW.d[27] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_00896_),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\dpath.RF.R[12][11] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_01581_),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\dpath.RF.R[18][30] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_00636_),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\dpath.RF.R[18][19] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_00625_),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\dpath.RF.R[22][25] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_00375_),
    .X(net1373));
 sky130_fd_sc_hd__buf_1 hold479 (.A(\dpath.RF.wdata[2] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_01212_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_00739_),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\dpath.RF.R[10][27] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_00860_),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\dpath.RF.R[9][4] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_00709_),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\dpath.RF.R[2][25] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_00826_),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\dpath.RF.R[28][30] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_00895_),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\dpath.RF.R[18][29] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\ctrl.inst_M[20] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_00635_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\dpath.RF.R[26][22] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_00919_),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\dpath.RF.R[22][28] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_00378_),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\dpath.RF.R[21][8] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_00422_),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\dpath.RF.R[21][1] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_00415_),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\dpath.RF.R[16][9] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\dpath.csrw_out_DX.q[31] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_00306_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_00551_),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\dpath.RF.R[18][22] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_00628_),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\dpath.RF.R[20][5] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_00483_),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\dpath.RF.R[1][10] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_00520_),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\dpath.RF.R[2][22] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_00823_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\dpath.RF.R[20][1] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\dpath.csrw_out_MW.d[6] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_00479_),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\dpath.RF.R[30][19] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_01658_),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\dpath.RF.R[26][29] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_00926_),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\dpath.RF.R[22][20] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_00370_),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\dpath.RF.R[19][2] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_00320_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\dpath.RF.R[24][7] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_01191_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_01609_),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\dpath.RF.R[10][4] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_00837_),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\dpath.RF.R[14][26] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_01307_),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\dpath.RF.R[16][2] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_00544_),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\dpath.RF.R[14][8] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_01289_),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\dpath.RF.R[1][0] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\dpath.csrw_out_DX.q[21] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_00510_),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\dpath.RF.R[1][29] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_00539_),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\dpath.RF.R[17][20] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_00466_),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\dpath.RF.R[14][31] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_01312_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\dpath.RF.R[1][19] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_00529_),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\dpath.RF.R[16][16] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_01462_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_00558_),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\dpath.RF.R[2][18] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_00819_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\dpath.RF.R[26][7] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_00904_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\dpath.RF.R[17][16] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_00462_),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\dpath.RF.R[18][25] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_00631_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\dpath.RF.R[9][19] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\dpath.csrw_out_MW.d[7] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_00724_),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\dpath.RF.R[12][22] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_01592_),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\dpath.RF.R[14][27] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_01308_),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\dpath.RF.R[22][12] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_00362_),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\dpath.RF.R[2][31] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_00832_),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\dpath.RF.R[1][22] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_01192_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_00532_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\dpath.RF.R[19][10] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_00328_),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\dpath.RF.R[8][27] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_01020_),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\dpath.RF.R[6][19] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_00061_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\dpath.RF.R[17][25] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_00471_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\dpath.RF.R[10][9] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\dpath.csrw_out_DX.q[22] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_00842_),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\dpath.RF.R[26][31] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_00928_),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\ctrl.inst_X[6] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_00242_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\dpath.RF.R[30][28] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_01667_),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\dpath.RF.R[21][9] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_00423_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\dpath.RF.R[26][9] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_01463_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_00906_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\dpath.RF.R[12][14] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_01584_),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\dpath.RF.R[18][18] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_00624_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\dpath.RF.R[2][16] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_00817_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\dpath.RF.R[23][18] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_00686_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\dpath.RF.R[8][0] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\dpath.csrw_out_DX.q[20] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_00993_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\dpath.RF.R[18][0] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_00606_),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\dpath.RF.R[20][22] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_00500_),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\dpath.RF.R[16][3] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_00545_),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\dpath.RF.R[28][13] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_00878_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\dpath.RF.R[20][28] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_01472_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_01461_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_00506_),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\dpath.RF.R[17][15] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_00461_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\dpath.RF.R[16][4] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_00546_),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\dpath.RF.R[22][15] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_00365_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\dpath.RF.R[28][23] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_00888_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\dpath.RF.R[24][15] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\dpath.csrw_out_MW.d[3] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_01617_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\dpath.RF.R[20][12] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_00490_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\dpath.RF.R[2][19] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_00820_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\dpath.RF.R[10][20] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_00853_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\dpath.RF.R[5][20] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_00222_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\dpath.RF.R[20][0] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_01188_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_00478_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\dpath.RF.R[5][21] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_00223_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\dpath.RF.R[2][27] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_00828_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\dpath.RF.R[13][24] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_01497_),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\dpath.RF.R[1][25] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_00535_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\dpath.RF.R[16][29] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\dpath.csrw_out_MW.d[0] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_00571_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\dpath.RF.R[16][11] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_00553_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\dpath.RF.R[22][27] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_00377_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\dpath.RF.R[30][2] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_01641_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\dpath.RF.R[1][17] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_00527_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\dpath.RF.R[8][14] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_01185_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_01007_),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\dpath.RF.R[24][6] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_01608_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\dpath.RF.R[18][20] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_00626_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\dpath.RF.R[22][23] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_00373_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\dpath.RF.R[12][7] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_01577_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\dpath.RF.R[9][23] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\ctrl.inst_M[31] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_00728_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\dpath.RF.R[28][28] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_00893_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\dpath.RF.R[25][14] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_00751_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\dpath.RF.R[26][30] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_00927_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\dpath.RF.R[16][30] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_00572_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\dpath.RF.R[6][20] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_00317_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_00062_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\dpath.RF.R[30][5] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_01644_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\dpath.RF.R[6][18] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_00060_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\dpath.RF.R[8][9] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_01002_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\dpath.RF.R[17][28] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_00474_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\dpath.RF.R[9][15] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\dpath.csrw_out_MW.d[11] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_00720_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\dpath.RF.R[26][4] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_00901_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\dpath.RF.R[20][18] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_00496_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\dpath.RF.R[5][22] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_00224_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\dpath.RF.R[13][30] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_01503_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\dpath.RF.R[24][23] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_01196_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_01625_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\dpath.RF.R[5][3] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_00205_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\dpath.RF.R[9][26] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_00731_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\dpath.RF.R[6][23] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_00065_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\dpath.RF.R[6][11] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_00053_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\dpath.RF.R[14][18] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\dpath.csrw_out_MW.d[2] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_01299_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\dpath.RF.R[22][22] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_00372_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\dpath.RF.R[25][17] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_00754_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\dpath.RF.R[12][19] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_01589_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\dpath.RF.R[2][13] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_00814_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\dpath.RF.R[17][22] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\dpath.csrw_out_DX.q[8] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_01187_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_00468_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\dpath.RF.R[22][14] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_00364_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\dpath.RF.R[2][28] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_00829_),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\dpath.RF.R[13][11] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_01484_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\dpath.csrw_out_MW.d[31] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_01216_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\dpath.RF.R[9][8] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\dpath.csrw_out_MW.d[14] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_00713_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\dpath.RF.R[24][9] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_01611_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\dpath.RF.R[5][15] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_00217_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\dpath.RF.R[30][27] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_01666_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\dpath.RF.R[5][7] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_00209_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\dpath.RF.R[26][3] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_01199_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_00900_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\dpath.RF.R[28][19] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_00884_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\dpath.RF.R[30][17] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_01656_),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\dpath.RF.R[9][13] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_00718_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\dpath.RF.R[10][29] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_00862_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\dpath.RF.R[23][22] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\dpath.csrw_out_MW.d[15] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_00690_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\dpath.RF.R[26][28] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_00925_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\dpath.RF.R[17][8] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_00454_),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\dpath.RF.R[16][27] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_00569_),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\dpath.RF.R[26][15] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_00912_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\dpath.RF.R[6][25] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_01200_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_00067_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\dpath.RF.R[14][24] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_01305_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\dpath.RF.R[1][1] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_00511_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\dpath.RF.R[7][7] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_00017_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\dpath.RF.R[18][15] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_00621_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\dpath.RF.R[25][9] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\dpath.csrw_out_MW.d[17] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_00746_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\dpath.RF.R[22][4] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_00354_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\dpath.RF.R[14][29] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_01310_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\dpath.RF.R[6][1] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_00043_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\dpath.RF.R[20][15] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_00493_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\dpath.RF.R[19][27] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_01202_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_00345_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\dpath.RF.R[7][25] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_00035_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\dpath.RF.R[10][2] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_00835_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\dpath.RF.R[30][10] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_01649_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\dpath.RF.R[12][16] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_01586_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\dpath.RF.R[13][31] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\ctrl.inst_M[1] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_01504_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\dpath.RF.R[28][24] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_00889_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\dpath.RF.R[27][27] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_00988_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\dpath.RF.R[5][27] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_00229_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\dpath.RF.R[24][11] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_01613_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\dpath.RF.R[18][4] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_00292_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_00610_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\dpath.RF.R[18][11] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_00617_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\dpath.RF.R[24][30] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_01632_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\dpath.RF.R[8][13] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_01006_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\dpath.RF.R[10][31] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_00864_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\dpath.RF.R[9][5] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\dpath.csrw_out_MW.d[26] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_00710_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\dpath.RF.R[28][14] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_00879_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\dpath.RF.R[8][22] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_01015_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\dpath.RF.R[27][30] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_00991_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\dpath.RF.R[17][29] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_00475_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\dpath.RF.R[20][14] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_01449_),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_01211_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_00492_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\dpath.RF.R[21][7] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_00421_),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\dpath.RF.R[24][12] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_01614_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\dpath.RF.R[20][20] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_00498_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\dpath.RF.R[24][28] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_01630_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\dpath.RF.R[6][4] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\dpath.csrw_out_MW.d[10] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_00046_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\dpath.RF.R[30][4] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_01643_),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\dpath.RF.R[20][29] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_00507_),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\dpath.RF.R[26][8] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_00905_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\dpath.RF.R[1][11] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_00521_),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\dpath.RF.R[24][26] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_01195_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_01628_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\dpath.RF.R[20][10] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_00488_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\dpath.RF.R[21][30] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_00444_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\dpath.RF.R[22][29] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_00379_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\dpath.RF.R[25][26] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_00763_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\dpath.RF.R[30][29] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\dpath.csrw_out_MW.d[18] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_01668_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\dpath.RF.R[17][10] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_00456_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\dpath.RF.R[30][26] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_01665_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\dpath.RF.R[21][28] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_00442_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\dpath.RF.R[14][22] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_01303_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\dpath.RF.R[5][23] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_01203_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_00225_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\dpath.RF.R[18][23] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_00629_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\dpath.RF.R[12][24] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_01594_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\dpath.RF.R[12][15] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_01585_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\dpath.RF.R[10][23] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_00856_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\dpath.RF.R[9][27] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\dpath.csrw_out_DX.q[15] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_00732_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\dpath.RF.R[16][7] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_00549_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\dpath.RF.R[28][1] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_00866_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\dpath.RF.R[10][0] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_00833_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\dpath.RF.R[19][15] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_00333_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\dpath.RF.R[6][2] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_01456_),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_00044_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\dpath.RF.R[2][4] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_00805_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\dpath.RF.R[27][18] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_00979_),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\dpath.RF.R[11][21] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_00950_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\dpath.RF.R[7][23] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_00033_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\dpath.RF.R[25][27] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\dpath.csrw_out_MW.d[25] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_00764_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\dpath.RF.R[6][31] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_00073_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\dpath.RF.R[23][17] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_00685_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\dpath.RF.R[9][30] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_00735_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\dpath.RF.R[28][29] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_00894_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\dpath.RF.R[24][19] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_01210_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_01621_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\dpath.RF.R[30][15] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_01654_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\dpath.RF.R[12][1] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_01571_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\dpath.RF.R[18][31] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_00637_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\dpath.RF.R[10][14] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_00847_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\dpath.RF.R[14][9] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\dpath.csrw_out_DX.q[18] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_01290_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\dpath.RF.R[5][11] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_00213_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\dpath.RF.R[12][5] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_01575_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\dpath.RF.R[19][1] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_00319_),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\dpath.RF.R[18][24] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_00630_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\dpath.RF.R[22][10] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\dpath.csrw_out_DX.q[17] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_01459_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_00360_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\dpath.RF.R[25][7] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_00744_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\dpath.RF.R[17][27] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_00473_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\dpath.RF.R[6][8] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_00050_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\dpath.RF.R[2][1] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_00802_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\dpath.RF.R[24][14] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\dpath.sd_DX.q[7] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_01616_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\dpath.RF.R[26][18] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_00915_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\dpath.RF.R[17][6] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_00452_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\dpath.RF.R[30][20] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_01659_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\dpath.RF.R[12][0] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_01570_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\dpath.RF.R[10][24] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_00389_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_00857_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\dpath.RF.R[28][21] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_00886_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\dpath.RF.R[10][3] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_00836_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\dpath.RF.R[18][9] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_00615_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\dpath.RF.R[14][13] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_01294_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\dpath.RF.R[7][4] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\dpath.csrw_out_MW.d[21] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_00014_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\dpath.RF.R[16][22] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_00564_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\dpath.RF.R[26][20] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_00917_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\dpath.RF.R[14][3] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_01284_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\dpath.RF.R[8][15] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_01008_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\dpath.RF.R[9][3] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_01206_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_00708_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\dpath.RF.R[19][20] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_00338_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\dpath.RF.R[14][16] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_01297_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\dpath.RF.R[6][29] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_00071_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\dpath.RF.R[13][15] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_01488_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\dpath.RF.R[12][4] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\ctrl.inst_X[26] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_01574_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\dpath.RF.R[13][22] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_01495_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\dpath.RF.R[12][30] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_01600_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\dpath.RF.R[30][12] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_01651_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\dpath.RF.R[28][3] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_00868_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\dpath.RF.R[18][10] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_00257_),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_00616_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\dpath.RF.R[1][26] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_00536_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\dpath.RF.R[13][28] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_01501_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\dpath.RF.R[28][10] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_00875_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\dpath.RF.R[11][10] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_00939_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\dpath.RF.R[18][13] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\dpath.csrw_out_DX.q[14] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_00619_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\dpath.RF.R[2][3] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_00804_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\dpath.RF.R[17][11] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_00457_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\dpath.RF.R[29][2] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_00140_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\dpath.RF.R[18][17] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_00623_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\dpath.RF.R[20][21] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_01455_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_00499_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\dpath.RF.R[14][11] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_01292_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\dpath.RF.R[25][25] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_00762_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\dpath.RF.R[19][0] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_00318_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\dpath.RF.R[26][16] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_00913_),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\dpath.RF.R[16][13] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\dpath.csrw_out_DX.q[26] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_00555_),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\dpath.RF.R[11][31] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_00960_),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\dpath.RF.R[20][11] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_00489_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\dpath.RF.R[10][6] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_00839_),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\dpath.RF.R[28][12] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_00877_),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\dpath.RF.R[23][28] ),
    .X(net1894));
 sky130_fd_sc_hd__buf_2 input1 (.A(dmemresp_rdata[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(dmemresp_rdata[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(in1[12]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(in1[13]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(in1[14]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(in1[15]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(in1[16]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(in1[17]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(in1[18]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(in1[19]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(in1[1]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(in1[20]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(dmemresp_rdata[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(in1[21]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(in1[22]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(in1[23]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(in1[24]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(in1[25]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(in1[26]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(in1[27]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(in1[28]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(in1[29]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(in1[2]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(dmemresp_rdata[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(in1[30]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(in1[31]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(in1[3]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(in1[4]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(in1[5]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(in1[6]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(in1[7]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(in1[8]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(in1[9]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(in2[0]),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(dmemresp_rdata[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(in2[10]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(in2[11]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(in2[12]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(in2[13]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(in2[14]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(in2[15]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(in2[16]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(in2[17]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(in2[18]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(in2[19]),
    .X(net139));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(dmemresp_rdata[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(in2[1]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(in2[20]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(in2[21]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(in2[22]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(in2[23]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(in2[24]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(in2[25]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(in2[26]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(in2[27]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(in2[28]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(dmemresp_rdata[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(in2[29]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 input151 (.A(in2[2]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(in2[30]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 input153 (.A(in2[31]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(in2[3]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 input155 (.A(in2[4]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(in2[5]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 input157 (.A(in2[6]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 input158 (.A(in2[7]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(in2[8]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(dmemresp_rdata[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(in2[9]),
    .X(net160));
 sky130_fd_sc_hd__dlymetal6s2s_1 input161 (.A(rst),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(dmemresp_rdata[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(dmemresp_rdata[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(dmemresp_rdata[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(dmemresp_rdata[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(dmemresp_rdata[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(dmemresp_rdata[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(dmemresp_rdata[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(dmemresp_rdata[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(dmemresp_rdata[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(dmemresp_rdata[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(dmemresp_rdata[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(dmemresp_rdata[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(dmemresp_rdata[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(dmemresp_rdata[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(dmemresp_rdata[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(dmemresp_rdata[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(dmemresp_rdata[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(dmemresp_rdata[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(imemresp_data[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(imemresp_data[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(imemresp_data[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(imemresp_data[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(imemresp_data[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(imemresp_data[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(imemresp_data[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(dmemresp_rdata[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(imemresp_data[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(imemresp_data[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(imemresp_data[18]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(imemresp_data[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(imemresp_data[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(imemresp_data[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(imemresp_data[21]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(imemresp_data[22]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(imemresp_data[23]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(imemresp_data[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(dmemresp_rdata[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(imemresp_data[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(imemresp_data[26]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(imemresp_data[27]),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 input53 (.A(imemresp_data[28]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(imemresp_data[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(imemresp_data[2]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(imemresp_data[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(imemresp_data[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(imemresp_data[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(imemresp_data[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(dmemresp_rdata[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(imemresp_data[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(imemresp_data[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(imemresp_data[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(imemresp_data[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(imemresp_data[9]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(in0[0]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(in0[10]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(in0[11]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(in0[12]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(in0[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(dmemresp_rdata[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input70 (.A(in0[14]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(in0[15]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(in0[16]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(in0[17]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(in0[18]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(in0[19]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(in0[1]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(in0[20]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(in0[21]),
    .X(net78));
 sky130_fd_sc_hd__dlymetal6s2s_1 input79 (.A(in0[22]),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(dmemresp_rdata[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input80 (.A(in0[23]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(in0[24]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(in0[25]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(in0[26]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(in0[27]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(in0[28]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(in0[29]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(in0[2]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(in0[30]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(in0[31]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(dmemresp_rdata[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input90 (.A(in0[3]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(in0[4]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(in0[5]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(in0[6]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(in0[7]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(in0[8]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(in0[9]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(in1[0]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(in1[10]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(in1[11]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 max_cap356 (.A(_05453_),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 max_cap481 (.A(_01971_),
    .X(net481));
 sky130_fd_sc_hd__buf_4 max_cap486 (.A(_02070_),
    .X(net486));
 sky130_fd_sc_hd__buf_12 output162 (.A(net162),
    .X(dmemreq_addr[0]));
 sky130_fd_sc_hd__buf_12 output163 (.A(net163),
    .X(dmemreq_addr[10]));
 sky130_fd_sc_hd__buf_12 output164 (.A(net164),
    .X(dmemreq_addr[11]));
 sky130_fd_sc_hd__buf_12 output165 (.A(net165),
    .X(dmemreq_addr[12]));
 sky130_fd_sc_hd__buf_12 output166 (.A(net166),
    .X(dmemreq_addr[13]));
 sky130_fd_sc_hd__buf_12 output167 (.A(net167),
    .X(dmemreq_addr[14]));
 sky130_fd_sc_hd__buf_12 output168 (.A(net168),
    .X(dmemreq_addr[15]));
 sky130_fd_sc_hd__buf_12 output169 (.A(net169),
    .X(dmemreq_addr[16]));
 sky130_fd_sc_hd__buf_12 output170 (.A(net170),
    .X(dmemreq_addr[17]));
 sky130_fd_sc_hd__buf_12 output171 (.A(net171),
    .X(dmemreq_addr[18]));
 sky130_fd_sc_hd__buf_12 output172 (.A(net172),
    .X(dmemreq_addr[19]));
 sky130_fd_sc_hd__buf_12 output173 (.A(net173),
    .X(dmemreq_addr[1]));
 sky130_fd_sc_hd__buf_12 output174 (.A(net174),
    .X(dmemreq_addr[20]));
 sky130_fd_sc_hd__buf_12 output175 (.A(net175),
    .X(dmemreq_addr[21]));
 sky130_fd_sc_hd__buf_12 output176 (.A(net176),
    .X(dmemreq_addr[22]));
 sky130_fd_sc_hd__buf_12 output177 (.A(net177),
    .X(dmemreq_addr[23]));
 sky130_fd_sc_hd__buf_12 output178 (.A(net178),
    .X(dmemreq_addr[24]));
 sky130_fd_sc_hd__buf_12 output179 (.A(net179),
    .X(dmemreq_addr[25]));
 sky130_fd_sc_hd__buf_12 output180 (.A(net180),
    .X(dmemreq_addr[26]));
 sky130_fd_sc_hd__buf_12 output181 (.A(net181),
    .X(dmemreq_addr[27]));
 sky130_fd_sc_hd__buf_12 output182 (.A(net182),
    .X(dmemreq_addr[28]));
 sky130_fd_sc_hd__buf_12 output183 (.A(net183),
    .X(dmemreq_addr[29]));
 sky130_fd_sc_hd__buf_12 output184 (.A(net184),
    .X(dmemreq_addr[2]));
 sky130_fd_sc_hd__buf_12 output185 (.A(net185),
    .X(dmemreq_addr[30]));
 sky130_fd_sc_hd__buf_12 output186 (.A(net186),
    .X(dmemreq_addr[31]));
 sky130_fd_sc_hd__buf_12 output187 (.A(net187),
    .X(dmemreq_addr[3]));
 sky130_fd_sc_hd__buf_12 output188 (.A(net188),
    .X(dmemreq_addr[4]));
 sky130_fd_sc_hd__buf_12 output189 (.A(net189),
    .X(dmemreq_addr[5]));
 sky130_fd_sc_hd__buf_12 output190 (.A(net190),
    .X(dmemreq_addr[6]));
 sky130_fd_sc_hd__buf_12 output191 (.A(net191),
    .X(dmemreq_addr[7]));
 sky130_fd_sc_hd__buf_12 output192 (.A(net192),
    .X(dmemreq_addr[8]));
 sky130_fd_sc_hd__buf_12 output193 (.A(net193),
    .X(dmemreq_addr[9]));
 sky130_fd_sc_hd__buf_12 output194 (.A(net194),
    .X(dmemreq_type));
 sky130_fd_sc_hd__buf_12 output195 (.A(net195),
    .X(dmemreq_val));
 sky130_fd_sc_hd__buf_12 output196 (.A(net196),
    .X(dmemreq_wdata[0]));
 sky130_fd_sc_hd__buf_12 output197 (.A(net197),
    .X(dmemreq_wdata[10]));
 sky130_fd_sc_hd__buf_12 output198 (.A(net198),
    .X(dmemreq_wdata[11]));
 sky130_fd_sc_hd__buf_12 output199 (.A(net199),
    .X(dmemreq_wdata[12]));
 sky130_fd_sc_hd__buf_12 output200 (.A(net200),
    .X(dmemreq_wdata[13]));
 sky130_fd_sc_hd__buf_12 output201 (.A(net201),
    .X(dmemreq_wdata[14]));
 sky130_fd_sc_hd__buf_12 output202 (.A(net202),
    .X(dmemreq_wdata[15]));
 sky130_fd_sc_hd__buf_12 output203 (.A(net203),
    .X(dmemreq_wdata[16]));
 sky130_fd_sc_hd__buf_12 output204 (.A(net204),
    .X(dmemreq_wdata[17]));
 sky130_fd_sc_hd__buf_12 output205 (.A(net205),
    .X(dmemreq_wdata[18]));
 sky130_fd_sc_hd__buf_12 output206 (.A(net206),
    .X(dmemreq_wdata[19]));
 sky130_fd_sc_hd__buf_12 output207 (.A(net207),
    .X(dmemreq_wdata[1]));
 sky130_fd_sc_hd__buf_12 output208 (.A(net208),
    .X(dmemreq_wdata[20]));
 sky130_fd_sc_hd__buf_12 output209 (.A(net209),
    .X(dmemreq_wdata[21]));
 sky130_fd_sc_hd__buf_12 output210 (.A(net210),
    .X(dmemreq_wdata[22]));
 sky130_fd_sc_hd__buf_12 output211 (.A(net211),
    .X(dmemreq_wdata[23]));
 sky130_fd_sc_hd__buf_12 output212 (.A(net212),
    .X(dmemreq_wdata[24]));
 sky130_fd_sc_hd__buf_12 output213 (.A(net213),
    .X(dmemreq_wdata[25]));
 sky130_fd_sc_hd__buf_12 output214 (.A(net214),
    .X(dmemreq_wdata[26]));
 sky130_fd_sc_hd__buf_12 output215 (.A(net215),
    .X(dmemreq_wdata[27]));
 sky130_fd_sc_hd__buf_12 output216 (.A(net216),
    .X(dmemreq_wdata[28]));
 sky130_fd_sc_hd__buf_12 output217 (.A(net217),
    .X(dmemreq_wdata[29]));
 sky130_fd_sc_hd__buf_12 output218 (.A(net218),
    .X(dmemreq_wdata[2]));
 sky130_fd_sc_hd__buf_12 output219 (.A(net219),
    .X(dmemreq_wdata[30]));
 sky130_fd_sc_hd__buf_12 output220 (.A(net220),
    .X(dmemreq_wdata[31]));
 sky130_fd_sc_hd__buf_12 output221 (.A(net221),
    .X(dmemreq_wdata[3]));
 sky130_fd_sc_hd__buf_12 output222 (.A(net222),
    .X(dmemreq_wdata[4]));
 sky130_fd_sc_hd__buf_12 output223 (.A(net223),
    .X(dmemreq_wdata[5]));
 sky130_fd_sc_hd__buf_12 output224 (.A(net224),
    .X(dmemreq_wdata[6]));
 sky130_fd_sc_hd__buf_12 output225 (.A(net225),
    .X(dmemreq_wdata[7]));
 sky130_fd_sc_hd__buf_12 output226 (.A(net226),
    .X(dmemreq_wdata[8]));
 sky130_fd_sc_hd__buf_12 output227 (.A(net227),
    .X(dmemreq_wdata[9]));
 sky130_fd_sc_hd__buf_12 output228 (.A(net228),
    .X(imemreq_addr[0]));
 sky130_fd_sc_hd__buf_12 output229 (.A(net229),
    .X(imemreq_addr[10]));
 sky130_fd_sc_hd__buf_12 output230 (.A(net230),
    .X(imemreq_addr[11]));
 sky130_fd_sc_hd__buf_12 output231 (.A(net231),
    .X(imemreq_addr[12]));
 sky130_fd_sc_hd__buf_12 output232 (.A(net232),
    .X(imemreq_addr[13]));
 sky130_fd_sc_hd__buf_12 output233 (.A(net233),
    .X(imemreq_addr[14]));
 sky130_fd_sc_hd__buf_12 output234 (.A(net234),
    .X(imemreq_addr[15]));
 sky130_fd_sc_hd__buf_12 output235 (.A(net235),
    .X(imemreq_addr[16]));
 sky130_fd_sc_hd__buf_12 output236 (.A(net236),
    .X(imemreq_addr[17]));
 sky130_fd_sc_hd__buf_12 output237 (.A(net237),
    .X(imemreq_addr[18]));
 sky130_fd_sc_hd__buf_12 output238 (.A(net238),
    .X(imemreq_addr[19]));
 sky130_fd_sc_hd__buf_12 output239 (.A(net239),
    .X(imemreq_addr[1]));
 sky130_fd_sc_hd__buf_12 output240 (.A(net240),
    .X(imemreq_addr[20]));
 sky130_fd_sc_hd__buf_12 output241 (.A(net241),
    .X(imemreq_addr[21]));
 sky130_fd_sc_hd__buf_12 output242 (.A(net242),
    .X(imemreq_addr[22]));
 sky130_fd_sc_hd__buf_12 output243 (.A(net243),
    .X(imemreq_addr[23]));
 sky130_fd_sc_hd__buf_12 output244 (.A(net244),
    .X(imemreq_addr[24]));
 sky130_fd_sc_hd__buf_12 output245 (.A(net245),
    .X(imemreq_addr[25]));
 sky130_fd_sc_hd__buf_12 output246 (.A(net246),
    .X(imemreq_addr[26]));
 sky130_fd_sc_hd__buf_12 output247 (.A(net247),
    .X(imemreq_addr[27]));
 sky130_fd_sc_hd__buf_12 output248 (.A(net248),
    .X(imemreq_addr[28]));
 sky130_fd_sc_hd__buf_12 output249 (.A(net249),
    .X(imemreq_addr[29]));
 sky130_fd_sc_hd__buf_12 output250 (.A(net250),
    .X(imemreq_addr[2]));
 sky130_fd_sc_hd__buf_12 output251 (.A(net251),
    .X(imemreq_addr[30]));
 sky130_fd_sc_hd__buf_12 output252 (.A(net252),
    .X(imemreq_addr[31]));
 sky130_fd_sc_hd__buf_12 output253 (.A(net253),
    .X(imemreq_addr[3]));
 sky130_fd_sc_hd__buf_12 output254 (.A(net254),
    .X(imemreq_addr[4]));
 sky130_fd_sc_hd__buf_12 output255 (.A(net255),
    .X(imemreq_addr[5]));
 sky130_fd_sc_hd__buf_12 output256 (.A(net256),
    .X(imemreq_addr[6]));
 sky130_fd_sc_hd__buf_12 output257 (.A(net257),
    .X(imemreq_addr[7]));
 sky130_fd_sc_hd__buf_12 output258 (.A(net258),
    .X(imemreq_addr[8]));
 sky130_fd_sc_hd__buf_12 output259 (.A(net259),
    .X(imemreq_addr[9]));
 sky130_fd_sc_hd__buf_12 output260 (.A(net260),
    .X(out0[0]));
 sky130_fd_sc_hd__buf_12 output261 (.A(net261),
    .X(out0[10]));
 sky130_fd_sc_hd__buf_12 output262 (.A(net262),
    .X(out0[11]));
 sky130_fd_sc_hd__buf_12 output263 (.A(net263),
    .X(out0[12]));
 sky130_fd_sc_hd__buf_12 output264 (.A(net264),
    .X(out0[13]));
 sky130_fd_sc_hd__buf_12 output265 (.A(net265),
    .X(out0[14]));
 sky130_fd_sc_hd__buf_12 output266 (.A(net266),
    .X(out0[15]));
 sky130_fd_sc_hd__buf_12 output267 (.A(net267),
    .X(out0[16]));
 sky130_fd_sc_hd__buf_12 output268 (.A(net268),
    .X(out0[17]));
 sky130_fd_sc_hd__buf_12 output269 (.A(net269),
    .X(out0[18]));
 sky130_fd_sc_hd__buf_12 output270 (.A(net270),
    .X(out0[19]));
 sky130_fd_sc_hd__buf_12 output271 (.A(net271),
    .X(out0[1]));
 sky130_fd_sc_hd__buf_12 output272 (.A(net272),
    .X(out0[20]));
 sky130_fd_sc_hd__buf_12 output273 (.A(net273),
    .X(out0[21]));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(out0[22]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(out0[23]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(out0[24]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(out0[25]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(out0[26]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(out0[27]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(out0[28]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(out0[29]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(out0[2]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(out0[30]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(out0[31]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(out0[3]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(out0[4]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(out0[5]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(out0[6]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(out0[7]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(out0[8]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(out0[9]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(out1[0]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(out1[10]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(out1[11]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(out1[12]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(out1[13]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(out1[14]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(out1[15]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(out1[16]));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(out1[17]));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(out1[18]));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(out1[19]));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(out1[1]));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(out1[20]));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(out1[21]));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(out1[22]));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(out1[23]));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(out1[24]));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(out1[25]));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(out1[26]));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(out1[27]));
 sky130_fd_sc_hd__buf_12 output312 (.A(net312),
    .X(out1[28]));
 sky130_fd_sc_hd__buf_12 output313 (.A(net313),
    .X(out1[29]));
 sky130_fd_sc_hd__buf_12 output314 (.A(net314),
    .X(out1[2]));
 sky130_fd_sc_hd__buf_12 output315 (.A(net315),
    .X(out1[30]));
 sky130_fd_sc_hd__buf_12 output316 (.A(net316),
    .X(out1[31]));
 sky130_fd_sc_hd__buf_12 output317 (.A(net317),
    .X(out1[3]));
 sky130_fd_sc_hd__buf_12 output318 (.A(net318),
    .X(out1[4]));
 sky130_fd_sc_hd__buf_12 output319 (.A(net319),
    .X(out1[5]));
 sky130_fd_sc_hd__buf_12 output320 (.A(net320),
    .X(out1[6]));
 sky130_fd_sc_hd__buf_12 output321 (.A(net321),
    .X(out1[7]));
 sky130_fd_sc_hd__buf_12 output322 (.A(net322),
    .X(out1[8]));
 sky130_fd_sc_hd__buf_12 output323 (.A(net323),
    .X(out1[9]));
 sky130_fd_sc_hd__buf_12 output324 (.A(net324),
    .X(out2[0]));
 sky130_fd_sc_hd__buf_12 output325 (.A(net325),
    .X(out2[10]));
 sky130_fd_sc_hd__buf_12 output326 (.A(net326),
    .X(out2[11]));
 sky130_fd_sc_hd__buf_12 output327 (.A(net327),
    .X(out2[12]));
 sky130_fd_sc_hd__buf_12 output328 (.A(net328),
    .X(out2[13]));
 sky130_fd_sc_hd__buf_12 output329 (.A(net329),
    .X(out2[14]));
 sky130_fd_sc_hd__buf_12 output330 (.A(net330),
    .X(out2[15]));
 sky130_fd_sc_hd__buf_12 output331 (.A(net331),
    .X(out2[16]));
 sky130_fd_sc_hd__buf_12 output332 (.A(net332),
    .X(out2[17]));
 sky130_fd_sc_hd__buf_12 output333 (.A(net333),
    .X(out2[18]));
 sky130_fd_sc_hd__buf_12 output334 (.A(net334),
    .X(out2[19]));
 sky130_fd_sc_hd__buf_12 output335 (.A(net335),
    .X(out2[1]));
 sky130_fd_sc_hd__buf_12 output336 (.A(net336),
    .X(out2[20]));
 sky130_fd_sc_hd__buf_12 output337 (.A(net337),
    .X(out2[21]));
 sky130_fd_sc_hd__buf_12 output338 (.A(net338),
    .X(out2[22]));
 sky130_fd_sc_hd__buf_12 output339 (.A(net339),
    .X(out2[23]));
 sky130_fd_sc_hd__buf_12 output340 (.A(net340),
    .X(out2[24]));
 sky130_fd_sc_hd__buf_12 output341 (.A(net341),
    .X(out2[25]));
 sky130_fd_sc_hd__buf_12 output342 (.A(net342),
    .X(out2[26]));
 sky130_fd_sc_hd__buf_12 output343 (.A(net343),
    .X(out2[27]));
 sky130_fd_sc_hd__buf_12 output344 (.A(net344),
    .X(out2[28]));
 sky130_fd_sc_hd__buf_12 output345 (.A(net345),
    .X(out2[29]));
 sky130_fd_sc_hd__buf_12 output346 (.A(net346),
    .X(out2[2]));
 sky130_fd_sc_hd__buf_12 output347 (.A(net347),
    .X(out2[30]));
 sky130_fd_sc_hd__buf_12 output348 (.A(net348),
    .X(out2[31]));
 sky130_fd_sc_hd__buf_12 output349 (.A(net349),
    .X(out2[3]));
 sky130_fd_sc_hd__buf_12 output350 (.A(net350),
    .X(out2[4]));
 sky130_fd_sc_hd__buf_12 output351 (.A(net351),
    .X(out2[5]));
 sky130_fd_sc_hd__buf_12 output352 (.A(net352),
    .X(out2[6]));
 sky130_fd_sc_hd__buf_12 output353 (.A(net353),
    .X(out2[7]));
 sky130_fd_sc_hd__buf_12 output354 (.A(net354),
    .X(out2[8]));
 sky130_fd_sc_hd__buf_12 output355 (.A(net355),
    .X(out2[9]));
 assign imemreq_val = net895;
endmodule

